
// 	Wed May  5 22:49:17 2021
//	vlsi
//	localhost.localdomain

module Pooling_2x2_Routing (start, \image_in[0][0] , \image_in[0][1] , \image_in[0][2] , 
    \image_in[0][3] , \image_in[0][4] , \image_in[1][0] , \image_in[1][1] , \image_in[1][2] , 
    \image_in[1][3] , \image_in[1][4] , \image_in[2][0] , \image_in[2][1] , \image_in[2][2] , 
    \image_in[2][3] , \image_in[2][4] , \image_in[3][0] , \image_in[3][1] , \image_in[3][2] , 
    \image_in[3][3] , \image_in[3][4] , \image_in[4][0] , \image_in[4][1] , \image_in[4][2] , 
    \image_in[4][3] , \image_in[4][4] , finish, pixel_out);

output finish;
output [15:0] pixel_out;
input [15:0] \image_in[0][0] ;
input [15:0] \image_in[0][1] ;
input [15:0] \image_in[0][2] ;
input [15:0] \image_in[0][3] ;
input [15:0] \image_in[0][4] ;
input [15:0] \image_in[1][0] ;
input [15:0] \image_in[1][1] ;
input [15:0] \image_in[1][2] ;
input [15:0] \image_in[1][3] ;
input [15:0] \image_in[1][4] ;
input [15:0] \image_in[2][0] ;
input [15:0] \image_in[2][1] ;
input [15:0] \image_in[2][2] ;
input [15:0] \image_in[2][3] ;
input [15:0] \image_in[2][4] ;
input [15:0] \image_in[3][0] ;
input [15:0] \image_in[3][1] ;
input [15:0] \image_in[3][2] ;
input [15:0] \image_in[3][3] ;
input [15:0] \image_in[3][4] ;
input [15:0] \image_in[4][0] ;
input [15:0] \image_in[4][1] ;
input [15:0] \image_in[4][2] ;
input [15:0] \image_in[4][3] ;
input [15:0] \image_in[4][4] ;
input start;
wire n_0_0_0;
wire n_0_0_1;
wire n_0_0_2;
wire n_0_0_3;
wire n_0_0_4;
wire n_0_0_5;
wire n_0_0_6;
wire n_0_0_7;
wire n_0_0_8;
wire n_0_0_9;
wire n_0_0_10;
wire n_0_0_11;
wire n_0_0_12;
wire n_0_0_13;
wire n_0_0_14;
wire n_0_0_15;
wire n_0_0_16;
wire n_0_0_17;
wire n_0_0_18;
wire n_0_0_19;
wire n_0_0_20;
wire n_0_0_21;
wire n_0_0_22;
wire n_0_0_23;
wire n_0_0_24;
wire n_0_0_25;
wire n_0_0_26;
wire n_0_0_27;
wire n_0_0_28;
wire n_0_0_29;
wire n_0_0_30;
wire n_0_0_31;
wire n_0_0_32;
wire n_0_0_33;
wire n_0_0_34;
wire n_0_0_35;
wire n_0_0_36;
wire n_0_0_37;
wire n_0_0_38;
wire n_0_0_39;
wire n_0_0_40;
wire n_0_0_41;
wire n_0_0_42;
wire n_0_0_43;
wire n_0_0_44;
wire n_0_0_45;
wire n_0_0_46;
wire n_0_0_47;
wire n_0_0_48;
wire n_0_0_49;
wire n_0_0_50;
wire n_0_0_51;
wire n_0_0_52;
wire n_0_0_53;
wire n_0_0_54;
wire n_0_0_55;
wire n_0_0_56;
wire n_0_0_57;
wire n_0_0_62;
wire n_0_0_63;
wire n_0_0_64;
wire n_0_0_65;
wire n_0_0_58;
wire n_0_0_66;
wire n_0_0_59;
wire n_0_0_67;
wire n_0_0_60;
wire n_0_0_68;
wire n_0_0_61;
wire n_0_0_69;
wire n_0_0_79;
wire n_0_0_70;
wire n_0_0_80;
wire n_0_0_71;
wire n_0_0_81;
wire n_0_0_72;
wire n_0_0_82;
wire n_0_0_73;
wire n_0_0_83;
wire n_0_0_74;
wire n_0_0_84;
wire n_0_0_75;
wire n_0_0_85;
wire n_0_0_76;
wire n_0_0_86;
wire n_0_0_77;
wire n_0_0_87;
wire n_0_0_78;
wire n_0_0_88;
wire n_0_0_89;
wire n_0_0_90;
wire n_0_0_91;
wire n_0_0_92;
wire n_0_0_93;

assign finish = start;
// WARNING . Detected multiport output net(s). Introducing ASSIGN statements.
// This may cause simulation/synthesis mismatches . 
assign pixel_out[15] = 1'b0 ;
assign pixel_out[14] = 1'b0 ;

XNOR2_X1 i_0_0_63 (.ZN (n_0_0_93), .A (\image_in[1][0] [15] ), .B (\image_in[1][1] [15] ));
XNOR2_X1 i_0_0_62 (.ZN (n_0_0_92), .A (n_0_0_57), .B (n_0_0_78));
XNOR2_X1 i_0_0_61 (.ZN (n_0_0_91), .A (n_0_0_93), .B (n_0_0_92));
XOR2_X1 i_0_0_60 (.Z (n_0_0_90), .A (\image_in[0][0] [15] ), .B (n_0_0_55));
XNOR2_X1 i_0_0_59 (.ZN (n_0_0_89), .A (\image_in[0][1] [15] ), .B (n_0_0_90));
OAI21_X1 i_0_0_58 (.ZN (n_0_0_88), .A (start), .B1 (n_0_0_91), .B2 (n_0_0_89));
AOI21_X1 i_0_0_57 (.ZN (pixel_out[13]), .A (n_0_0_88), .B1 (n_0_0_89), .B2 (n_0_0_91));
AND2_X1 i_0_0_56 (.ZN (pixel_out[12]), .A1 (start), .A2 (n_0_0_87));
AND2_X1 i_0_0_55 (.ZN (pixel_out[11]), .A1 (start), .A2 (n_0_0_86));
AND2_X1 i_0_0_54 (.ZN (pixel_out[10]), .A1 (start), .A2 (n_0_0_85));
AND2_X1 i_0_0_53 (.ZN (pixel_out[9]), .A1 (start), .A2 (n_0_0_84));
AND2_X1 i_0_0_52 (.ZN (pixel_out[8]), .A1 (start), .A2 (n_0_0_83));
AND2_X1 i_0_0_51 (.ZN (pixel_out[7]), .A1 (start), .A2 (n_0_0_82));
AND2_X1 i_0_0_50 (.ZN (pixel_out[6]), .A1 (start), .A2 (n_0_0_81));
AND2_X1 i_0_0_49 (.ZN (pixel_out[5]), .A1 (start), .A2 (n_0_0_80));
AND2_X1 i_0_0_48 (.ZN (pixel_out[4]), .A1 (start), .A2 (n_0_0_79));
AND2_X1 i_0_0_47 (.ZN (pixel_out[3]), .A1 (start), .A2 (n_0_0_61));
AND2_X1 i_0_0_46 (.ZN (pixel_out[2]), .A1 (start), .A2 (n_0_0_60));
AND2_X1 i_0_0_45 (.ZN (pixel_out[1]), .A1 (start), .A2 (n_0_0_59));
AND2_X1 i_0_0_44 (.ZN (pixel_out[0]), .A1 (start), .A2 (n_0_0_58));
FA_X1 i_0_0_43 (.CO (n_0_0_78), .S (n_0_0_87), .A (n_0_0_53), .B (n_0_0_56), .CI (n_0_0_77));
FA_X1 i_0_0_42 (.CO (n_0_0_77), .S (n_0_0_86), .A (n_0_0_49), .B (n_0_0_52), .CI (n_0_0_76));
FA_X1 i_0_0_41 (.CO (n_0_0_76), .S (n_0_0_85), .A (n_0_0_45), .B (n_0_0_48), .CI (n_0_0_75));
FA_X1 i_0_0_40 (.CO (n_0_0_75), .S (n_0_0_84), .A (n_0_0_41), .B (n_0_0_44), .CI (n_0_0_74));
FA_X1 i_0_0_39 (.CO (n_0_0_74), .S (n_0_0_83), .A (n_0_0_37), .B (n_0_0_40), .CI (n_0_0_73));
FA_X1 i_0_0_38 (.CO (n_0_0_73), .S (n_0_0_82), .A (n_0_0_33), .B (n_0_0_36), .CI (n_0_0_72));
FA_X1 i_0_0_37 (.CO (n_0_0_72), .S (n_0_0_81), .A (n_0_0_29), .B (n_0_0_32), .CI (n_0_0_71));
FA_X1 i_0_0_36 (.CO (n_0_0_71), .S (n_0_0_80), .A (n_0_0_25), .B (n_0_0_28), .CI (n_0_0_70));
FA_X1 i_0_0_35 (.CO (n_0_0_70), .S (n_0_0_79), .A (n_0_0_21), .B (n_0_0_24), .CI (n_0_0_69));
FA_X1 i_0_0_34 (.CO (n_0_0_69), .S (n_0_0_61), .A (n_0_0_17), .B (n_0_0_20), .CI (n_0_0_68));
FA_X1 i_0_0_33 (.CO (n_0_0_68), .S (n_0_0_60), .A (n_0_0_13), .B (n_0_0_16), .CI (n_0_0_67));
FA_X1 i_0_0_32 (.CO (n_0_0_67), .S (n_0_0_59), .A (n_0_0_10), .B (n_0_0_12), .CI (n_0_0_66));
FA_X1 i_0_0_31 (.CO (n_0_0_66), .S (n_0_0_58), .A (n_0_0_6), .B (n_0_0_8), .CI (n_0_0_65));
FA_X1 i_0_0_30 (.CO (n_0_0_65), .S (n_0_0_64), .A (n_0_0_4), .B (n_0_0_2), .CI (n_0_0_63));
HA_X1 i_0_0_29 (.CO (n_0_0_63), .S (n_0_0_62), .A (\image_in[0][0] [0] ), .B (n_0_0_0));
FA_X1 i_0_0_28 (.CO (n_0_0_57), .S (n_0_0_56), .A (\image_in[0][0] [14] ), .B (n_0_0_51), .CI (n_0_0_54));
FA_X1 i_0_0_27 (.CO (n_0_0_55), .S (n_0_0_54), .A (\image_in[0][1] [14] ), .B (\image_in[1][0] [14] ), .CI (\image_in[1][1] [14] ));
FA_X1 i_0_0_26 (.CO (n_0_0_53), .S (n_0_0_52), .A (\image_in[0][0] [13] ), .B (n_0_0_47), .CI (n_0_0_50));
FA_X1 i_0_0_25 (.CO (n_0_0_51), .S (n_0_0_50), .A (\image_in[0][1] [13] ), .B (\image_in[1][0] [13] ), .CI (\image_in[1][1] [13] ));
FA_X1 i_0_0_24 (.CO (n_0_0_49), .S (n_0_0_48), .A (\image_in[0][0] [12] ), .B (n_0_0_43), .CI (n_0_0_46));
FA_X1 i_0_0_23 (.CO (n_0_0_47), .S (n_0_0_46), .A (\image_in[0][1] [12] ), .B (\image_in[1][0] [12] ), .CI (\image_in[1][1] [12] ));
FA_X1 i_0_0_22 (.CO (n_0_0_45), .S (n_0_0_44), .A (\image_in[0][0] [11] ), .B (n_0_0_39), .CI (n_0_0_42));
FA_X1 i_0_0_21 (.CO (n_0_0_43), .S (n_0_0_42), .A (\image_in[0][1] [11] ), .B (\image_in[1][0] [11] ), .CI (\image_in[1][1] [11] ));
FA_X1 i_0_0_20 (.CO (n_0_0_41), .S (n_0_0_40), .A (\image_in[0][0] [10] ), .B (n_0_0_35), .CI (n_0_0_38));
FA_X1 i_0_0_19 (.CO (n_0_0_39), .S (n_0_0_38), .A (\image_in[0][1] [10] ), .B (\image_in[1][0] [10] ), .CI (\image_in[1][1] [10] ));
FA_X1 i_0_0_18 (.CO (n_0_0_37), .S (n_0_0_36), .A (\image_in[0][0] [9] ), .B (n_0_0_31), .CI (n_0_0_34));
FA_X1 i_0_0_17 (.CO (n_0_0_35), .S (n_0_0_34), .A (\image_in[0][1] [9] ), .B (\image_in[1][0] [9] ), .CI (\image_in[1][1] [9] ));
FA_X1 i_0_0_16 (.CO (n_0_0_33), .S (n_0_0_32), .A (\image_in[0][0] [8] ), .B (n_0_0_27), .CI (n_0_0_30));
FA_X1 i_0_0_15 (.CO (n_0_0_31), .S (n_0_0_30), .A (\image_in[0][1] [8] ), .B (\image_in[1][0] [8] ), .CI (\image_in[1][1] [8] ));
FA_X1 i_0_0_14 (.CO (n_0_0_29), .S (n_0_0_28), .A (\image_in[0][0] [7] ), .B (n_0_0_23), .CI (n_0_0_26));
FA_X1 i_0_0_13 (.CO (n_0_0_27), .S (n_0_0_26), .A (\image_in[0][1] [7] ), .B (\image_in[1][0] [7] ), .CI (\image_in[1][1] [7] ));
FA_X1 i_0_0_12 (.CO (n_0_0_25), .S (n_0_0_24), .A (\image_in[0][0] [6] ), .B (n_0_0_19), .CI (n_0_0_22));
FA_X1 i_0_0_11 (.CO (n_0_0_23), .S (n_0_0_22), .A (\image_in[0][1] [6] ), .B (\image_in[1][0] [6] ), .CI (\image_in[1][1] [6] ));
FA_X1 i_0_0_10 (.CO (n_0_0_21), .S (n_0_0_20), .A (\image_in[0][0] [5] ), .B (n_0_0_15), .CI (n_0_0_18));
FA_X1 i_0_0_9 (.CO (n_0_0_19), .S (n_0_0_18), .A (\image_in[0][1] [5] ), .B (\image_in[1][0] [5] ), .CI (\image_in[1][1] [5] ));
FA_X1 i_0_0_8 (.CO (n_0_0_17), .S (n_0_0_16), .A (\image_in[0][0] [4] ), .B (n_0_0_11), .CI (n_0_0_14));
FA_X1 i_0_0_7 (.CO (n_0_0_15), .S (n_0_0_14), .A (\image_in[0][1] [4] ), .B (\image_in[1][0] [4] ), .CI (\image_in[1][1] [4] ));
FA_X1 i_0_0_6 (.CO (n_0_0_13), .S (n_0_0_12), .A (\image_in[0][0] [3] ), .B (n_0_0_7), .CI (n_0_0_9));
FA_X1 i_0_0_5 (.CO (n_0_0_11), .S (n_0_0_10), .A (\image_in[0][1] [3] ), .B (\image_in[1][0] [3] ), .CI (\image_in[1][1] [3] ));
FA_X1 i_0_0_4 (.CO (n_0_0_9), .S (n_0_0_8), .A (\image_in[0][0] [2] ), .B (n_0_0_3), .CI (n_0_0_5));
FA_X1 i_0_0_3 (.CO (n_0_0_7), .S (n_0_0_6), .A (\image_in[0][1] [2] ), .B (\image_in[1][0] [2] ), .CI (\image_in[1][1] [2] ));
HA_X1 i_0_0_2 (.CO (n_0_0_5), .S (n_0_0_4), .A (\image_in[0][0] [1] ), .B (n_0_0_1));
FA_X1 i_0_0_1 (.CO (n_0_0_3), .S (n_0_0_2), .A (\image_in[0][1] [1] ), .B (\image_in[1][0] [1] ), .CI (\image_in[1][1] [1] ));
FA_X1 i_0_0_0 (.CO (n_0_0_1), .S (n_0_0_0), .A (\image_in[0][1] [0] ), .B (\image_in[1][0] [0] ), .CI (\image_in[1][1] [0] ));

endmodule //Pooling_2x2


