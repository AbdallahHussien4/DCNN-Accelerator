/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Wed May  5 21:50:23 2021
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 1812433378 */

module datapath__0_2(p_0, p_1, p_2);
   input [32:0]p_0;
   input [32:0]p_1;
   output [32:0]p_2;

   HA_X1 i_1 (.A(p_0[17]), .B(p_1[17]), .CO(n_1), .S(p_2[17]));
   FA_X1 i_2 (.A(p_0[18]), .B(p_1[18]), .CI(n_1), .CO(n_2), .S(p_2[18]));
   FA_X1 i_3 (.A(p_0[19]), .B(p_1[19]), .CI(n_2), .CO(n_3), .S(p_2[19]));
   FA_X1 i_4 (.A(p_0[20]), .B(p_1[20]), .CI(n_3), .CO(n_4), .S(p_2[20]));
   FA_X1 i_5 (.A(p_0[21]), .B(p_1[21]), .CI(n_4), .CO(n_5), .S(p_2[21]));
   FA_X1 i_6 (.A(p_0[22]), .B(p_1[22]), .CI(n_5), .CO(n_6), .S(p_2[22]));
   FA_X1 i_7 (.A(p_0[23]), .B(p_1[23]), .CI(n_6), .CO(n_7), .S(p_2[23]));
   FA_X1 i_8 (.A(p_0[24]), .B(p_1[24]), .CI(n_7), .CO(n_8), .S(p_2[24]));
   FA_X1 i_9 (.A(p_0[25]), .B(p_1[25]), .CI(n_8), .CO(n_9), .S(p_2[25]));
   FA_X1 i_10 (.A(p_0[26]), .B(p_1[26]), .CI(n_9), .CO(n_10), .S(p_2[26]));
   FA_X1 i_11 (.A(p_0[27]), .B(p_1[27]), .CI(n_10), .CO(n_11), .S(p_2[27]));
   FA_X1 i_12 (.A(p_0[28]), .B(p_1[28]), .CI(n_11), .CO(n_12), .S(p_2[28]));
   FA_X1 i_13 (.A(p_0[29]), .B(p_1[29]), .CI(n_12), .CO(n_13), .S(p_2[29]));
   FA_X1 i_14 (.A(p_0[30]), .B(p_1[30]), .CI(n_13), .CO(n_14), .S(p_2[30]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[31]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[31]), .B1(p_0[31]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[32]), .B(n_15), .Z(p_2[32]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[31]), .A3(n_16), .B1(p_0[31]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[31]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[31]), .ZN(n_18));
endmodule

module datapath__0_3(p_0, p_1, p_2);
   input [32:0]p_0;
   input [32:0]p_1;
   output [32:0]p_2;

   HA_X1 i_1 (.A(p_0[17]), .B(p_1[17]), .CO(n_1), .S(p_2[17]));
   FA_X1 i_2 (.A(p_0[18]), .B(p_1[18]), .CI(n_1), .CO(n_2), .S(p_2[18]));
   FA_X1 i_3 (.A(p_0[19]), .B(p_1[19]), .CI(n_2), .CO(n_3), .S(p_2[19]));
   FA_X1 i_4 (.A(p_0[20]), .B(p_1[20]), .CI(n_3), .CO(n_4), .S(p_2[20]));
   FA_X1 i_5 (.A(p_0[21]), .B(p_1[21]), .CI(n_4), .CO(n_5), .S(p_2[21]));
   FA_X1 i_6 (.A(p_0[22]), .B(p_1[22]), .CI(n_5), .CO(n_6), .S(p_2[22]));
   FA_X1 i_7 (.A(p_0[23]), .B(p_1[23]), .CI(n_6), .CO(n_7), .S(p_2[23]));
   FA_X1 i_8 (.A(p_0[24]), .B(p_1[24]), .CI(n_7), .CO(n_8), .S(p_2[24]));
   FA_X1 i_9 (.A(p_0[25]), .B(p_1[25]), .CI(n_8), .CO(n_9), .S(p_2[25]));
   FA_X1 i_10 (.A(p_0[26]), .B(p_1[26]), .CI(n_9), .CO(n_10), .S(p_2[26]));
   FA_X1 i_11 (.A(p_0[27]), .B(p_1[27]), .CI(n_10), .CO(n_11), .S(p_2[27]));
   FA_X1 i_12 (.A(p_0[28]), .B(p_1[28]), .CI(n_11), .CO(n_12), .S(p_2[28]));
   FA_X1 i_13 (.A(p_0[29]), .B(p_1[29]), .CI(n_12), .CO(n_13), .S(p_2[29]));
   FA_X1 i_14 (.A(p_0[30]), .B(p_1[30]), .CI(n_13), .CO(n_14), .S(p_2[30]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[31]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[31]), .B1(p_0[31]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[32]), .B(n_15), .Z(p_2[32]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[31]), .A3(n_16), .B1(p_0[31]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[31]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[31]), .ZN(n_18));
endmodule

module datapath__0_6(p_0, p_1, p_2);
   input [32:0]p_0;
   input [32:0]p_1;
   output [32:0]p_2;

   HA_X1 i_1 (.A(p_0[17]), .B(p_1[17]), .CO(n_1), .S(p_2[17]));
   FA_X1 i_2 (.A(p_0[18]), .B(p_1[18]), .CI(n_1), .CO(n_2), .S(p_2[18]));
   FA_X1 i_3 (.A(p_0[19]), .B(p_1[19]), .CI(n_2), .CO(n_3), .S(p_2[19]));
   FA_X1 i_4 (.A(p_0[20]), .B(p_1[20]), .CI(n_3), .CO(n_4), .S(p_2[20]));
   FA_X1 i_5 (.A(p_0[21]), .B(p_1[21]), .CI(n_4), .CO(n_5), .S(p_2[21]));
   FA_X1 i_6 (.A(p_0[22]), .B(p_1[22]), .CI(n_5), .CO(n_6), .S(p_2[22]));
   FA_X1 i_7 (.A(p_0[23]), .B(p_1[23]), .CI(n_6), .CO(n_7), .S(p_2[23]));
   FA_X1 i_8 (.A(p_0[24]), .B(p_1[24]), .CI(n_7), .CO(n_8), .S(p_2[24]));
   FA_X1 i_9 (.A(p_0[25]), .B(p_1[25]), .CI(n_8), .CO(n_9), .S(p_2[25]));
   FA_X1 i_10 (.A(p_0[26]), .B(p_1[26]), .CI(n_9), .CO(n_10), .S(p_2[26]));
   FA_X1 i_11 (.A(p_0[27]), .B(p_1[27]), .CI(n_10), .CO(n_11), .S(p_2[27]));
   FA_X1 i_12 (.A(p_0[28]), .B(p_1[28]), .CI(n_11), .CO(n_12), .S(p_2[28]));
   FA_X1 i_13 (.A(p_0[29]), .B(p_1[29]), .CI(n_12), .CO(n_13), .S(p_2[29]));
   FA_X1 i_14 (.A(p_0[30]), .B(p_1[30]), .CI(n_13), .CO(n_14), .S(p_2[30]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[31]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[31]), .B1(p_0[31]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[32]), .B(n_15), .Z(p_2[32]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[31]), .A3(n_16), .B1(p_0[31]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[31]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[31]), .ZN(n_18));
endmodule

module datapath__0_7(p_0, p_1, p_2);
   input [32:0]p_0;
   input [32:0]p_1;
   output [32:0]p_2;

   HA_X1 i_1 (.A(p_0[17]), .B(p_1[17]), .CO(n_1), .S(p_2[17]));
   FA_X1 i_2 (.A(p_0[18]), .B(p_1[18]), .CI(n_1), .CO(n_2), .S(p_2[18]));
   FA_X1 i_3 (.A(p_0[19]), .B(p_1[19]), .CI(n_2), .CO(n_3), .S(p_2[19]));
   FA_X1 i_4 (.A(p_0[20]), .B(p_1[20]), .CI(n_3), .CO(n_4), .S(p_2[20]));
   FA_X1 i_5 (.A(p_0[21]), .B(p_1[21]), .CI(n_4), .CO(n_5), .S(p_2[21]));
   FA_X1 i_6 (.A(p_0[22]), .B(p_1[22]), .CI(n_5), .CO(n_6), .S(p_2[22]));
   FA_X1 i_7 (.A(p_0[23]), .B(p_1[23]), .CI(n_6), .CO(n_7), .S(p_2[23]));
   FA_X1 i_8 (.A(p_0[24]), .B(p_1[24]), .CI(n_7), .CO(n_8), .S(p_2[24]));
   FA_X1 i_9 (.A(p_0[25]), .B(p_1[25]), .CI(n_8), .CO(n_9), .S(p_2[25]));
   FA_X1 i_10 (.A(p_0[26]), .B(p_1[26]), .CI(n_9), .CO(n_10), .S(p_2[26]));
   FA_X1 i_11 (.A(p_0[27]), .B(p_1[27]), .CI(n_10), .CO(n_11), .S(p_2[27]));
   FA_X1 i_12 (.A(p_0[28]), .B(p_1[28]), .CI(n_11), .CO(n_12), .S(p_2[28]));
   FA_X1 i_13 (.A(p_0[29]), .B(p_1[29]), .CI(n_12), .CO(n_13), .S(p_2[29]));
   FA_X1 i_14 (.A(p_0[30]), .B(p_1[30]), .CI(n_13), .CO(n_14), .S(p_2[30]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[31]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[31]), .B1(p_0[31]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[32]), .B(n_15), .Z(p_2[32]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[31]), .A3(n_16), .B1(p_0[31]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[31]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[31]), .ZN(n_18));
endmodule

module datapath__0_10(p_0, p_1, p_2);
   input [32:0]p_0;
   input [32:0]p_1;
   output [32:0]p_2;

   HA_X1 i_1 (.A(p_0[17]), .B(p_1[17]), .CO(n_1), .S(p_2[17]));
   FA_X1 i_2 (.A(p_0[18]), .B(p_1[18]), .CI(n_1), .CO(n_2), .S(p_2[18]));
   FA_X1 i_3 (.A(p_0[19]), .B(p_1[19]), .CI(n_2), .CO(n_3), .S(p_2[19]));
   FA_X1 i_4 (.A(p_0[20]), .B(p_1[20]), .CI(n_3), .CO(n_4), .S(p_2[20]));
   FA_X1 i_5 (.A(p_0[21]), .B(p_1[21]), .CI(n_4), .CO(n_5), .S(p_2[21]));
   FA_X1 i_6 (.A(p_0[22]), .B(p_1[22]), .CI(n_5), .CO(n_6), .S(p_2[22]));
   FA_X1 i_7 (.A(p_0[23]), .B(p_1[23]), .CI(n_6), .CO(n_7), .S(p_2[23]));
   FA_X1 i_8 (.A(p_0[24]), .B(p_1[24]), .CI(n_7), .CO(n_8), .S(p_2[24]));
   FA_X1 i_9 (.A(p_0[25]), .B(p_1[25]), .CI(n_8), .CO(n_9), .S(p_2[25]));
   FA_X1 i_10 (.A(p_0[26]), .B(p_1[26]), .CI(n_9), .CO(n_10), .S(p_2[26]));
   FA_X1 i_11 (.A(p_0[27]), .B(p_1[27]), .CI(n_10), .CO(n_11), .S(p_2[27]));
   FA_X1 i_12 (.A(p_0[28]), .B(p_1[28]), .CI(n_11), .CO(n_12), .S(p_2[28]));
   FA_X1 i_13 (.A(p_0[29]), .B(p_1[29]), .CI(n_12), .CO(n_13), .S(p_2[29]));
   FA_X1 i_14 (.A(p_0[30]), .B(p_1[30]), .CI(n_13), .CO(n_14), .S(p_2[30]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[31]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[31]), .B1(p_0[31]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[32]), .B(n_15), .Z(p_2[32]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[31]), .A3(n_16), .B1(p_0[31]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[31]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[31]), .ZN(n_18));
endmodule

module datapath__0_11(p_0, p_1, p_2);
   input [32:0]p_0;
   input [32:0]p_1;
   output [32:0]p_2;

   HA_X1 i_1 (.A(p_0[17]), .B(p_1[17]), .CO(n_1), .S(p_2[17]));
   FA_X1 i_2 (.A(p_0[18]), .B(p_1[18]), .CI(n_1), .CO(n_2), .S(p_2[18]));
   FA_X1 i_3 (.A(p_0[19]), .B(p_1[19]), .CI(n_2), .CO(n_3), .S(p_2[19]));
   FA_X1 i_4 (.A(p_0[20]), .B(p_1[20]), .CI(n_3), .CO(n_4), .S(p_2[20]));
   FA_X1 i_5 (.A(p_0[21]), .B(p_1[21]), .CI(n_4), .CO(n_5), .S(p_2[21]));
   FA_X1 i_6 (.A(p_0[22]), .B(p_1[22]), .CI(n_5), .CO(n_6), .S(p_2[22]));
   FA_X1 i_7 (.A(p_0[23]), .B(p_1[23]), .CI(n_6), .CO(n_7), .S(p_2[23]));
   FA_X1 i_8 (.A(p_0[24]), .B(p_1[24]), .CI(n_7), .CO(n_8), .S(p_2[24]));
   FA_X1 i_9 (.A(p_0[25]), .B(p_1[25]), .CI(n_8), .CO(n_9), .S(p_2[25]));
   FA_X1 i_10 (.A(p_0[26]), .B(p_1[26]), .CI(n_9), .CO(n_10), .S(p_2[26]));
   FA_X1 i_11 (.A(p_0[27]), .B(p_1[27]), .CI(n_10), .CO(n_11), .S(p_2[27]));
   FA_X1 i_12 (.A(p_0[28]), .B(p_1[28]), .CI(n_11), .CO(n_12), .S(p_2[28]));
   FA_X1 i_13 (.A(p_0[29]), .B(p_1[29]), .CI(n_12), .CO(n_13), .S(p_2[29]));
   FA_X1 i_14 (.A(p_0[30]), .B(p_1[30]), .CI(n_13), .CO(n_14), .S(p_2[30]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[31]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[31]), .B1(p_0[31]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[32]), .B(n_15), .Z(p_2[32]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[31]), .A3(n_16), .B1(p_0[31]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[31]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[31]), .ZN(n_18));
endmodule

module datapath__0_14(p_0, p_1, p_2);
   input [32:0]p_0;
   input [32:0]p_1;
   output [32:0]p_2;

   HA_X1 i_1 (.A(p_0[17]), .B(p_1[17]), .CO(n_1), .S(p_2[17]));
   FA_X1 i_2 (.A(p_0[18]), .B(p_1[18]), .CI(n_1), .CO(n_2), .S(p_2[18]));
   FA_X1 i_3 (.A(p_0[19]), .B(p_1[19]), .CI(n_2), .CO(n_3), .S(p_2[19]));
   FA_X1 i_4 (.A(p_0[20]), .B(p_1[20]), .CI(n_3), .CO(n_4), .S(p_2[20]));
   FA_X1 i_5 (.A(p_0[21]), .B(p_1[21]), .CI(n_4), .CO(n_5), .S(p_2[21]));
   FA_X1 i_6 (.A(p_0[22]), .B(p_1[22]), .CI(n_5), .CO(n_6), .S(p_2[22]));
   FA_X1 i_7 (.A(p_0[23]), .B(p_1[23]), .CI(n_6), .CO(n_7), .S(p_2[23]));
   FA_X1 i_8 (.A(p_0[24]), .B(p_1[24]), .CI(n_7), .CO(n_8), .S(p_2[24]));
   FA_X1 i_9 (.A(p_0[25]), .B(p_1[25]), .CI(n_8), .CO(n_9), .S(p_2[25]));
   FA_X1 i_10 (.A(p_0[26]), .B(p_1[26]), .CI(n_9), .CO(n_10), .S(p_2[26]));
   FA_X1 i_11 (.A(p_0[27]), .B(p_1[27]), .CI(n_10), .CO(n_11), .S(p_2[27]));
   FA_X1 i_12 (.A(p_0[28]), .B(p_1[28]), .CI(n_11), .CO(n_12), .S(p_2[28]));
   FA_X1 i_13 (.A(p_0[29]), .B(p_1[29]), .CI(n_12), .CO(n_13), .S(p_2[29]));
   FA_X1 i_14 (.A(p_0[30]), .B(p_1[30]), .CI(n_13), .CO(n_14), .S(p_2[30]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[31]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[31]), .B1(p_0[31]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[32]), .B(n_15), .Z(p_2[32]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[31]), .A3(n_16), .B1(p_0[31]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[31]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[31]), .ZN(n_18));
endmodule

module datapath__0_15(p_0, p_1, p_2);
   input [32:0]p_0;
   input [32:0]p_1;
   output [32:0]p_2;

   HA_X1 i_1 (.A(p_0[17]), .B(p_1[17]), .CO(n_1), .S(p_2[17]));
   FA_X1 i_2 (.A(p_0[18]), .B(p_1[18]), .CI(n_1), .CO(n_2), .S(p_2[18]));
   FA_X1 i_3 (.A(p_0[19]), .B(p_1[19]), .CI(n_2), .CO(n_3), .S(p_2[19]));
   FA_X1 i_4 (.A(p_0[20]), .B(p_1[20]), .CI(n_3), .CO(n_4), .S(p_2[20]));
   FA_X1 i_5 (.A(p_0[21]), .B(p_1[21]), .CI(n_4), .CO(n_5), .S(p_2[21]));
   FA_X1 i_6 (.A(p_0[22]), .B(p_1[22]), .CI(n_5), .CO(n_6), .S(p_2[22]));
   FA_X1 i_7 (.A(p_0[23]), .B(p_1[23]), .CI(n_6), .CO(n_7), .S(p_2[23]));
   FA_X1 i_8 (.A(p_0[24]), .B(p_1[24]), .CI(n_7), .CO(n_8), .S(p_2[24]));
   FA_X1 i_9 (.A(p_0[25]), .B(p_1[25]), .CI(n_8), .CO(n_9), .S(p_2[25]));
   FA_X1 i_10 (.A(p_0[26]), .B(p_1[26]), .CI(n_9), .CO(n_10), .S(p_2[26]));
   FA_X1 i_11 (.A(p_0[27]), .B(p_1[27]), .CI(n_10), .CO(n_11), .S(p_2[27]));
   FA_X1 i_12 (.A(p_0[28]), .B(p_1[28]), .CI(n_11), .CO(n_12), .S(p_2[28]));
   FA_X1 i_13 (.A(p_0[29]), .B(p_1[29]), .CI(n_12), .CO(n_13), .S(p_2[29]));
   FA_X1 i_14 (.A(p_0[30]), .B(p_1[30]), .CI(n_13), .CO(n_14), .S(p_2[30]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[31]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[31]), .B1(p_0[31]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[32]), .B(n_15), .Z(p_2[32]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[31]), .A3(n_16), .B1(p_0[31]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[31]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[31]), .ZN(n_18));
endmodule

module datapath__0_18(p_0, p_1, p_2);
   input [32:0]p_0;
   input [32:0]p_1;
   output [32:0]p_2;

   HA_X1 i_1 (.A(p_0[17]), .B(p_1[17]), .CO(n_1), .S(p_2[17]));
   FA_X1 i_2 (.A(p_0[18]), .B(p_1[18]), .CI(n_1), .CO(n_2), .S(p_2[18]));
   FA_X1 i_3 (.A(p_0[19]), .B(p_1[19]), .CI(n_2), .CO(n_3), .S(p_2[19]));
   FA_X1 i_4 (.A(p_0[20]), .B(p_1[20]), .CI(n_3), .CO(n_4), .S(p_2[20]));
   FA_X1 i_5 (.A(p_0[21]), .B(p_1[21]), .CI(n_4), .CO(n_5), .S(p_2[21]));
   FA_X1 i_6 (.A(p_0[22]), .B(p_1[22]), .CI(n_5), .CO(n_6), .S(p_2[22]));
   FA_X1 i_7 (.A(p_0[23]), .B(p_1[23]), .CI(n_6), .CO(n_7), .S(p_2[23]));
   FA_X1 i_8 (.A(p_0[24]), .B(p_1[24]), .CI(n_7), .CO(n_8), .S(p_2[24]));
   FA_X1 i_9 (.A(p_0[25]), .B(p_1[25]), .CI(n_8), .CO(n_9), .S(p_2[25]));
   FA_X1 i_10 (.A(p_0[26]), .B(p_1[26]), .CI(n_9), .CO(n_10), .S(p_2[26]));
   FA_X1 i_11 (.A(p_0[27]), .B(p_1[27]), .CI(n_10), .CO(n_11), .S(p_2[27]));
   FA_X1 i_12 (.A(p_0[28]), .B(p_1[28]), .CI(n_11), .CO(n_12), .S(p_2[28]));
   FA_X1 i_13 (.A(p_0[29]), .B(p_1[29]), .CI(n_12), .CO(n_13), .S(p_2[29]));
   FA_X1 i_14 (.A(p_0[30]), .B(p_1[30]), .CI(n_13), .CO(n_14), .S(p_2[30]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[31]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[31]), .B1(p_0[31]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[32]), .B(n_15), .Z(p_2[32]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[31]), .A3(n_16), .B1(p_0[31]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[31]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[31]), .ZN(n_18));
endmodule

module datapath__0_19(p_0, p_1, p_2);
   input [32:0]p_0;
   input [32:0]p_1;
   output [32:0]p_2;

   HA_X1 i_1 (.A(p_0[17]), .B(p_1[17]), .CO(n_1), .S(p_2[17]));
   FA_X1 i_2 (.A(p_0[18]), .B(p_1[18]), .CI(n_1), .CO(n_2), .S(p_2[18]));
   FA_X1 i_3 (.A(p_0[19]), .B(p_1[19]), .CI(n_2), .CO(n_3), .S(p_2[19]));
   FA_X1 i_4 (.A(p_0[20]), .B(p_1[20]), .CI(n_3), .CO(n_4), .S(p_2[20]));
   FA_X1 i_5 (.A(p_0[21]), .B(p_1[21]), .CI(n_4), .CO(n_5), .S(p_2[21]));
   FA_X1 i_6 (.A(p_0[22]), .B(p_1[22]), .CI(n_5), .CO(n_6), .S(p_2[22]));
   FA_X1 i_7 (.A(p_0[23]), .B(p_1[23]), .CI(n_6), .CO(n_7), .S(p_2[23]));
   FA_X1 i_8 (.A(p_0[24]), .B(p_1[24]), .CI(n_7), .CO(n_8), .S(p_2[24]));
   FA_X1 i_9 (.A(p_0[25]), .B(p_1[25]), .CI(n_8), .CO(n_9), .S(p_2[25]));
   FA_X1 i_10 (.A(p_0[26]), .B(p_1[26]), .CI(n_9), .CO(n_10), .S(p_2[26]));
   FA_X1 i_11 (.A(p_0[27]), .B(p_1[27]), .CI(n_10), .CO(n_11), .S(p_2[27]));
   FA_X1 i_12 (.A(p_0[28]), .B(p_1[28]), .CI(n_11), .CO(n_12), .S(p_2[28]));
   FA_X1 i_13 (.A(p_0[29]), .B(p_1[29]), .CI(n_12), .CO(n_13), .S(p_2[29]));
   FA_X1 i_14 (.A(p_0[30]), .B(p_1[30]), .CI(n_13), .CO(n_14), .S(p_2[30]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[31]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[31]), .B1(p_0[31]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[32]), .B(n_15), .Z(p_2[32]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[31]), .A3(n_16), .B1(p_0[31]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[31]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[31]), .ZN(n_18));
endmodule

module datapath__0_22(p_0, p_1, p_2);
   input [32:0]p_0;
   input [32:0]p_1;
   output [32:0]p_2;

   HA_X1 i_1 (.A(p_0[17]), .B(p_1[17]), .CO(n_1), .S(p_2[17]));
   FA_X1 i_2 (.A(p_0[18]), .B(p_1[18]), .CI(n_1), .CO(n_2), .S(p_2[18]));
   FA_X1 i_3 (.A(p_0[19]), .B(p_1[19]), .CI(n_2), .CO(n_3), .S(p_2[19]));
   FA_X1 i_4 (.A(p_0[20]), .B(p_1[20]), .CI(n_3), .CO(n_4), .S(p_2[20]));
   FA_X1 i_5 (.A(p_0[21]), .B(p_1[21]), .CI(n_4), .CO(n_5), .S(p_2[21]));
   FA_X1 i_6 (.A(p_0[22]), .B(p_1[22]), .CI(n_5), .CO(n_6), .S(p_2[22]));
   FA_X1 i_7 (.A(p_0[23]), .B(p_1[23]), .CI(n_6), .CO(n_7), .S(p_2[23]));
   FA_X1 i_8 (.A(p_0[24]), .B(p_1[24]), .CI(n_7), .CO(n_8), .S(p_2[24]));
   FA_X1 i_9 (.A(p_0[25]), .B(p_1[25]), .CI(n_8), .CO(n_9), .S(p_2[25]));
   FA_X1 i_10 (.A(p_0[26]), .B(p_1[26]), .CI(n_9), .CO(n_10), .S(p_2[26]));
   FA_X1 i_11 (.A(p_0[27]), .B(p_1[27]), .CI(n_10), .CO(n_11), .S(p_2[27]));
   FA_X1 i_12 (.A(p_0[28]), .B(p_1[28]), .CI(n_11), .CO(n_12), .S(p_2[28]));
   FA_X1 i_13 (.A(p_0[29]), .B(p_1[29]), .CI(n_12), .CO(n_13), .S(p_2[29]));
   FA_X1 i_14 (.A(p_0[30]), .B(p_1[30]), .CI(n_13), .CO(n_14), .S(p_2[30]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[31]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[31]), .B1(p_0[31]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[32]), .B(n_15), .Z(p_2[32]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[31]), .A3(n_16), .B1(p_0[31]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[31]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[31]), .ZN(n_18));
endmodule

module datapath__0_23(p_0, p_1, p_2);
   input [32:0]p_0;
   input [32:0]p_1;
   output [32:0]p_2;

   HA_X1 i_1 (.A(p_0[17]), .B(p_1[17]), .CO(n_1), .S(p_2[17]));
   FA_X1 i_2 (.A(p_0[18]), .B(p_1[18]), .CI(n_1), .CO(n_2), .S(p_2[18]));
   FA_X1 i_3 (.A(p_0[19]), .B(p_1[19]), .CI(n_2), .CO(n_3), .S(p_2[19]));
   FA_X1 i_4 (.A(p_0[20]), .B(p_1[20]), .CI(n_3), .CO(n_4), .S(p_2[20]));
   FA_X1 i_5 (.A(p_0[21]), .B(p_1[21]), .CI(n_4), .CO(n_5), .S(p_2[21]));
   FA_X1 i_6 (.A(p_0[22]), .B(p_1[22]), .CI(n_5), .CO(n_6), .S(p_2[22]));
   FA_X1 i_7 (.A(p_0[23]), .B(p_1[23]), .CI(n_6), .CO(n_7), .S(p_2[23]));
   FA_X1 i_8 (.A(p_0[24]), .B(p_1[24]), .CI(n_7), .CO(n_8), .S(p_2[24]));
   FA_X1 i_9 (.A(p_0[25]), .B(p_1[25]), .CI(n_8), .CO(n_9), .S(p_2[25]));
   FA_X1 i_10 (.A(p_0[26]), .B(p_1[26]), .CI(n_9), .CO(n_10), .S(p_2[26]));
   FA_X1 i_11 (.A(p_0[27]), .B(p_1[27]), .CI(n_10), .CO(n_11), .S(p_2[27]));
   FA_X1 i_12 (.A(p_0[28]), .B(p_1[28]), .CI(n_11), .CO(n_12), .S(p_2[28]));
   FA_X1 i_13 (.A(p_0[29]), .B(p_1[29]), .CI(n_12), .CO(n_13), .S(p_2[29]));
   FA_X1 i_14 (.A(p_0[30]), .B(p_1[30]), .CI(n_13), .CO(n_14), .S(p_2[30]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[31]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[31]), .B1(p_0[31]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[32]), .B(n_15), .Z(p_2[32]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[31]), .A3(n_16), .B1(p_0[31]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[31]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[31]), .ZN(n_18));
endmodule

module datapath__0_26(p_0, p_1, p_2);
   input [32:0]p_0;
   input [32:0]p_1;
   output [32:0]p_2;

   HA_X1 i_1 (.A(p_0[17]), .B(p_1[17]), .CO(n_1), .S(p_2[17]));
   FA_X1 i_2 (.A(p_0[18]), .B(p_1[18]), .CI(n_1), .CO(n_2), .S(p_2[18]));
   FA_X1 i_3 (.A(p_0[19]), .B(p_1[19]), .CI(n_2), .CO(n_3), .S(p_2[19]));
   FA_X1 i_4 (.A(p_0[20]), .B(p_1[20]), .CI(n_3), .CO(n_4), .S(p_2[20]));
   FA_X1 i_5 (.A(p_0[21]), .B(p_1[21]), .CI(n_4), .CO(n_5), .S(p_2[21]));
   FA_X1 i_6 (.A(p_0[22]), .B(p_1[22]), .CI(n_5), .CO(n_6), .S(p_2[22]));
   FA_X1 i_7 (.A(p_0[23]), .B(p_1[23]), .CI(n_6), .CO(n_7), .S(p_2[23]));
   FA_X1 i_8 (.A(p_0[24]), .B(p_1[24]), .CI(n_7), .CO(n_8), .S(p_2[24]));
   FA_X1 i_9 (.A(p_0[25]), .B(p_1[25]), .CI(n_8), .CO(n_9), .S(p_2[25]));
   FA_X1 i_10 (.A(p_0[26]), .B(p_1[26]), .CI(n_9), .CO(n_10), .S(p_2[26]));
   FA_X1 i_11 (.A(p_0[27]), .B(p_1[27]), .CI(n_10), .CO(n_11), .S(p_2[27]));
   FA_X1 i_12 (.A(p_0[28]), .B(p_1[28]), .CI(n_11), .CO(n_12), .S(p_2[28]));
   FA_X1 i_13 (.A(p_0[29]), .B(p_1[29]), .CI(n_12), .CO(n_13), .S(p_2[29]));
   FA_X1 i_14 (.A(p_0[30]), .B(p_1[30]), .CI(n_13), .CO(n_14), .S(p_2[30]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[31]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[31]), .B1(p_0[31]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[32]), .B(n_15), .Z(p_2[32]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[31]), .A3(n_16), .B1(p_0[31]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[31]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[31]), .ZN(n_18));
endmodule

module datapath__0_27(p_0, p_1, p_2);
   input [32:0]p_0;
   input [32:0]p_1;
   output [32:0]p_2;

   HA_X1 i_1 (.A(p_0[17]), .B(p_1[17]), .CO(n_1), .S(p_2[17]));
   FA_X1 i_2 (.A(p_0[18]), .B(p_1[18]), .CI(n_1), .CO(n_2), .S(p_2[18]));
   FA_X1 i_3 (.A(p_0[19]), .B(p_1[19]), .CI(n_2), .CO(n_3), .S(p_2[19]));
   FA_X1 i_4 (.A(p_0[20]), .B(p_1[20]), .CI(n_3), .CO(n_4), .S(p_2[20]));
   FA_X1 i_5 (.A(p_0[21]), .B(p_1[21]), .CI(n_4), .CO(n_5), .S(p_2[21]));
   FA_X1 i_6 (.A(p_0[22]), .B(p_1[22]), .CI(n_5), .CO(n_6), .S(p_2[22]));
   FA_X1 i_7 (.A(p_0[23]), .B(p_1[23]), .CI(n_6), .CO(n_7), .S(p_2[23]));
   FA_X1 i_8 (.A(p_0[24]), .B(p_1[24]), .CI(n_7), .CO(n_8), .S(p_2[24]));
   FA_X1 i_9 (.A(p_0[25]), .B(p_1[25]), .CI(n_8), .CO(n_9), .S(p_2[25]));
   FA_X1 i_10 (.A(p_0[26]), .B(p_1[26]), .CI(n_9), .CO(n_10), .S(p_2[26]));
   FA_X1 i_11 (.A(p_0[27]), .B(p_1[27]), .CI(n_10), .CO(n_11), .S(p_2[27]));
   FA_X1 i_12 (.A(p_0[28]), .B(p_1[28]), .CI(n_11), .CO(n_12), .S(p_2[28]));
   FA_X1 i_13 (.A(p_0[29]), .B(p_1[29]), .CI(n_12), .CO(n_13), .S(p_2[29]));
   FA_X1 i_14 (.A(p_0[30]), .B(p_1[30]), .CI(n_13), .CO(n_14), .S(p_2[30]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[31]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[31]), .B1(p_0[31]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[32]), .B(n_15), .Z(p_2[32]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[31]), .A3(n_16), .B1(p_0[31]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[31]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[31]), .ZN(n_18));
endmodule

module datapath__0_30(p_0, p_1, p_2);
   input [32:0]p_0;
   input [32:0]p_1;
   output [32:0]p_2;

   HA_X1 i_1 (.A(p_0[17]), .B(p_1[17]), .CO(n_1), .S(p_2[17]));
   FA_X1 i_2 (.A(p_0[18]), .B(p_1[18]), .CI(n_1), .CO(n_2), .S(p_2[18]));
   FA_X1 i_3 (.A(p_0[19]), .B(p_1[19]), .CI(n_2), .CO(n_3), .S(p_2[19]));
   FA_X1 i_4 (.A(p_0[20]), .B(p_1[20]), .CI(n_3), .CO(n_4), .S(p_2[20]));
   FA_X1 i_5 (.A(p_0[21]), .B(p_1[21]), .CI(n_4), .CO(n_5), .S(p_2[21]));
   FA_X1 i_6 (.A(p_0[22]), .B(p_1[22]), .CI(n_5), .CO(n_6), .S(p_2[22]));
   FA_X1 i_7 (.A(p_0[23]), .B(p_1[23]), .CI(n_6), .CO(n_7), .S(p_2[23]));
   FA_X1 i_8 (.A(p_0[24]), .B(p_1[24]), .CI(n_7), .CO(n_8), .S(p_2[24]));
   FA_X1 i_9 (.A(p_0[25]), .B(p_1[25]), .CI(n_8), .CO(n_9), .S(p_2[25]));
   FA_X1 i_10 (.A(p_0[26]), .B(p_1[26]), .CI(n_9), .CO(n_10), .S(p_2[26]));
   FA_X1 i_11 (.A(p_0[27]), .B(p_1[27]), .CI(n_10), .CO(n_11), .S(p_2[27]));
   FA_X1 i_12 (.A(p_0[28]), .B(p_1[28]), .CI(n_11), .CO(n_12), .S(p_2[28]));
   FA_X1 i_13 (.A(p_0[29]), .B(p_1[29]), .CI(n_12), .CO(n_13), .S(p_2[29]));
   FA_X1 i_14 (.A(p_0[30]), .B(p_1[30]), .CI(n_13), .CO(n_14), .S(p_2[30]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[31]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[31]), .B1(p_0[31]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[32]), .B(n_15), .Z(p_2[32]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[31]), .A3(n_16), .B1(p_0[31]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[31]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[31]), .ZN(n_18));
endmodule

module datapath__0_31(p_0, p_1, p_2);
   input [32:0]p_0;
   input [32:0]p_1;
   output [32:0]p_2;

   HA_X1 i_1 (.A(p_0[17]), .B(p_1[17]), .CO(n_1), .S(p_2[17]));
   FA_X1 i_2 (.A(p_0[18]), .B(p_1[18]), .CI(n_1), .CO(n_2), .S(p_2[18]));
   FA_X1 i_3 (.A(p_0[19]), .B(p_1[19]), .CI(n_2), .CO(n_3), .S(p_2[19]));
   FA_X1 i_4 (.A(p_0[20]), .B(p_1[20]), .CI(n_3), .CO(n_4), .S(p_2[20]));
   FA_X1 i_5 (.A(p_0[21]), .B(p_1[21]), .CI(n_4), .CO(n_5), .S(p_2[21]));
   FA_X1 i_6 (.A(p_0[22]), .B(p_1[22]), .CI(n_5), .CO(n_6), .S(p_2[22]));
   FA_X1 i_7 (.A(p_0[23]), .B(p_1[23]), .CI(n_6), .CO(n_7), .S(p_2[23]));
   FA_X1 i_8 (.A(p_0[24]), .B(p_1[24]), .CI(n_7), .CO(n_8), .S(p_2[24]));
   FA_X1 i_9 (.A(p_0[25]), .B(p_1[25]), .CI(n_8), .CO(n_9), .S(p_2[25]));
   FA_X1 i_10 (.A(p_0[26]), .B(p_1[26]), .CI(n_9), .CO(n_10), .S(p_2[26]));
   FA_X1 i_11 (.A(p_0[27]), .B(p_1[27]), .CI(n_10), .CO(n_11), .S(p_2[27]));
   FA_X1 i_12 (.A(p_0[28]), .B(p_1[28]), .CI(n_11), .CO(n_12), .S(p_2[28]));
   FA_X1 i_13 (.A(p_0[29]), .B(p_1[29]), .CI(n_12), .CO(n_13), .S(p_2[29]));
   FA_X1 i_14 (.A(p_0[30]), .B(p_1[30]), .CI(n_13), .CO(n_14), .S(p_2[30]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[31]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[31]), .B1(p_0[31]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[32]), .B(n_15), .Z(p_2[32]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[31]), .A3(n_16), .B1(p_0[31]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[31]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[31]), .ZN(n_18));
endmodule

module datapath__0_34(p_0, p_1, p_2);
   input [32:0]p_0;
   input [32:0]p_1;
   output [32:0]p_2;

   HA_X1 i_1 (.A(p_0[17]), .B(p_1[17]), .CO(n_1), .S(p_2[17]));
   FA_X1 i_2 (.A(p_0[18]), .B(p_1[18]), .CI(n_1), .CO(n_2), .S(p_2[18]));
   FA_X1 i_3 (.A(p_0[19]), .B(p_1[19]), .CI(n_2), .CO(n_3), .S(p_2[19]));
   FA_X1 i_4 (.A(p_0[20]), .B(p_1[20]), .CI(n_3), .CO(n_4), .S(p_2[20]));
   FA_X1 i_5 (.A(p_0[21]), .B(p_1[21]), .CI(n_4), .CO(n_5), .S(p_2[21]));
   FA_X1 i_6 (.A(p_0[22]), .B(p_1[22]), .CI(n_5), .CO(n_6), .S(p_2[22]));
   FA_X1 i_7 (.A(p_0[23]), .B(p_1[23]), .CI(n_6), .CO(n_7), .S(p_2[23]));
   FA_X1 i_8 (.A(p_0[24]), .B(p_1[24]), .CI(n_7), .CO(n_8), .S(p_2[24]));
   FA_X1 i_9 (.A(p_0[25]), .B(p_1[25]), .CI(n_8), .CO(n_9), .S(p_2[25]));
   FA_X1 i_10 (.A(p_0[26]), .B(p_1[26]), .CI(n_9), .CO(n_10), .S(p_2[26]));
   FA_X1 i_11 (.A(p_0[27]), .B(p_1[27]), .CI(n_10), .CO(n_11), .S(p_2[27]));
   FA_X1 i_12 (.A(p_0[28]), .B(p_1[28]), .CI(n_11), .CO(n_12), .S(p_2[28]));
   FA_X1 i_13 (.A(p_0[29]), .B(p_1[29]), .CI(n_12), .CO(n_13), .S(p_2[29]));
   FA_X1 i_14 (.A(p_0[30]), .B(p_1[30]), .CI(n_13), .CO(n_14), .S(p_2[30]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[31]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[31]), .B1(p_0[31]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[32]), .B(n_15), .Z(p_2[32]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[31]), .A3(n_16), .B1(p_0[31]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[31]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[31]), .ZN(n_18));
endmodule

module datapath__0_35(p_0, p_1, p_2);
   input [32:0]p_0;
   input [32:0]p_1;
   output [32:0]p_2;

   HA_X1 i_1 (.A(p_0[17]), .B(p_1[17]), .CO(n_1), .S(p_2[17]));
   FA_X1 i_2 (.A(p_0[18]), .B(p_1[18]), .CI(n_1), .CO(n_2), .S(p_2[18]));
   FA_X1 i_3 (.A(p_0[19]), .B(p_1[19]), .CI(n_2), .CO(n_3), .S(p_2[19]));
   FA_X1 i_4 (.A(p_0[20]), .B(p_1[20]), .CI(n_3), .CO(n_4), .S(p_2[20]));
   FA_X1 i_5 (.A(p_0[21]), .B(p_1[21]), .CI(n_4), .CO(n_5), .S(p_2[21]));
   FA_X1 i_6 (.A(p_0[22]), .B(p_1[22]), .CI(n_5), .CO(n_6), .S(p_2[22]));
   FA_X1 i_7 (.A(p_0[23]), .B(p_1[23]), .CI(n_6), .CO(n_7), .S(p_2[23]));
   FA_X1 i_8 (.A(p_0[24]), .B(p_1[24]), .CI(n_7), .CO(n_8), .S(p_2[24]));
   FA_X1 i_9 (.A(p_0[25]), .B(p_1[25]), .CI(n_8), .CO(n_9), .S(p_2[25]));
   FA_X1 i_10 (.A(p_0[26]), .B(p_1[26]), .CI(n_9), .CO(n_10), .S(p_2[26]));
   FA_X1 i_11 (.A(p_0[27]), .B(p_1[27]), .CI(n_10), .CO(n_11), .S(p_2[27]));
   FA_X1 i_12 (.A(p_0[28]), .B(p_1[28]), .CI(n_11), .CO(n_12), .S(p_2[28]));
   FA_X1 i_13 (.A(p_0[29]), .B(p_1[29]), .CI(n_12), .CO(n_13), .S(p_2[29]));
   FA_X1 i_14 (.A(p_0[30]), .B(p_1[30]), .CI(n_13), .CO(n_14), .S(p_2[30]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[31]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[31]), .B1(p_0[31]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[32]), .B(n_15), .Z(p_2[32]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[31]), .A3(n_16), .B1(p_0[31]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[31]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[31]), .ZN(n_18));
endmodule

module datapath__0_38(p_0, p_1, p_2);
   input [32:0]p_0;
   input [32:0]p_1;
   output [32:0]p_2;

   HA_X1 i_1 (.A(p_0[17]), .B(p_1[17]), .CO(n_1), .S(p_2[17]));
   FA_X1 i_2 (.A(p_0[18]), .B(p_1[18]), .CI(n_1), .CO(n_2), .S(p_2[18]));
   FA_X1 i_3 (.A(p_0[19]), .B(p_1[19]), .CI(n_2), .CO(n_3), .S(p_2[19]));
   FA_X1 i_4 (.A(p_0[20]), .B(p_1[20]), .CI(n_3), .CO(n_4), .S(p_2[20]));
   FA_X1 i_5 (.A(p_0[21]), .B(p_1[21]), .CI(n_4), .CO(n_5), .S(p_2[21]));
   FA_X1 i_6 (.A(p_0[22]), .B(p_1[22]), .CI(n_5), .CO(n_6), .S(p_2[22]));
   FA_X1 i_7 (.A(p_0[23]), .B(p_1[23]), .CI(n_6), .CO(n_7), .S(p_2[23]));
   FA_X1 i_8 (.A(p_0[24]), .B(p_1[24]), .CI(n_7), .CO(n_8), .S(p_2[24]));
   FA_X1 i_9 (.A(p_0[25]), .B(p_1[25]), .CI(n_8), .CO(n_9), .S(p_2[25]));
   FA_X1 i_10 (.A(p_0[26]), .B(p_1[26]), .CI(n_9), .CO(n_10), .S(p_2[26]));
   FA_X1 i_11 (.A(p_0[27]), .B(p_1[27]), .CI(n_10), .CO(n_11), .S(p_2[27]));
   FA_X1 i_12 (.A(p_0[28]), .B(p_1[28]), .CI(n_11), .CO(n_12), .S(p_2[28]));
   FA_X1 i_13 (.A(p_0[29]), .B(p_1[29]), .CI(n_12), .CO(n_13), .S(p_2[29]));
   FA_X1 i_14 (.A(p_0[30]), .B(p_1[30]), .CI(n_13), .CO(n_14), .S(p_2[30]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[31]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[31]), .B1(p_0[31]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[32]), .B(n_15), .Z(p_2[32]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[31]), .A3(n_16), .B1(p_0[31]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[31]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[31]), .ZN(n_18));
endmodule

module datapath__0_39(p_0, p_1, p_2);
   input [32:0]p_0;
   input [32:0]p_1;
   output [32:0]p_2;

   HA_X1 i_1 (.A(p_0[17]), .B(p_1[17]), .CO(n_1), .S(p_2[17]));
   FA_X1 i_2 (.A(p_0[18]), .B(p_1[18]), .CI(n_1), .CO(n_2), .S(p_2[18]));
   FA_X1 i_3 (.A(p_0[19]), .B(p_1[19]), .CI(n_2), .CO(n_3), .S(p_2[19]));
   FA_X1 i_4 (.A(p_0[20]), .B(p_1[20]), .CI(n_3), .CO(n_4), .S(p_2[20]));
   FA_X1 i_5 (.A(p_0[21]), .B(p_1[21]), .CI(n_4), .CO(n_5), .S(p_2[21]));
   FA_X1 i_6 (.A(p_0[22]), .B(p_1[22]), .CI(n_5), .CO(n_6), .S(p_2[22]));
   FA_X1 i_7 (.A(p_0[23]), .B(p_1[23]), .CI(n_6), .CO(n_7), .S(p_2[23]));
   FA_X1 i_8 (.A(p_0[24]), .B(p_1[24]), .CI(n_7), .CO(n_8), .S(p_2[24]));
   FA_X1 i_9 (.A(p_0[25]), .B(p_1[25]), .CI(n_8), .CO(n_9), .S(p_2[25]));
   FA_X1 i_10 (.A(p_0[26]), .B(p_1[26]), .CI(n_9), .CO(n_10), .S(p_2[26]));
   FA_X1 i_11 (.A(p_0[27]), .B(p_1[27]), .CI(n_10), .CO(n_11), .S(p_2[27]));
   FA_X1 i_12 (.A(p_0[28]), .B(p_1[28]), .CI(n_11), .CO(n_12), .S(p_2[28]));
   FA_X1 i_13 (.A(p_0[29]), .B(p_1[29]), .CI(n_12), .CO(n_13), .S(p_2[29]));
   FA_X1 i_14 (.A(p_0[30]), .B(p_1[30]), .CI(n_13), .CO(n_14), .S(p_2[30]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[31]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[31]), .B1(p_0[31]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[32]), .B(n_15), .Z(p_2[32]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[31]), .A3(n_16), .B1(p_0[31]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[31]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[31]), .ZN(n_18));
endmodule

module datapath__0_42(p_0, p_1, p_2);
   input [32:0]p_0;
   input [32:0]p_1;
   output [32:0]p_2;

   HA_X1 i_1 (.A(p_0[17]), .B(p_1[17]), .CO(n_1), .S(p_2[17]));
   FA_X1 i_2 (.A(p_0[18]), .B(p_1[18]), .CI(n_1), .CO(n_2), .S(p_2[18]));
   FA_X1 i_3 (.A(p_0[19]), .B(p_1[19]), .CI(n_2), .CO(n_3), .S(p_2[19]));
   FA_X1 i_4 (.A(p_0[20]), .B(p_1[20]), .CI(n_3), .CO(n_4), .S(p_2[20]));
   FA_X1 i_5 (.A(p_0[21]), .B(p_1[21]), .CI(n_4), .CO(n_5), .S(p_2[21]));
   FA_X1 i_6 (.A(p_0[22]), .B(p_1[22]), .CI(n_5), .CO(n_6), .S(p_2[22]));
   FA_X1 i_7 (.A(p_0[23]), .B(p_1[23]), .CI(n_6), .CO(n_7), .S(p_2[23]));
   FA_X1 i_8 (.A(p_0[24]), .B(p_1[24]), .CI(n_7), .CO(n_8), .S(p_2[24]));
   FA_X1 i_9 (.A(p_0[25]), .B(p_1[25]), .CI(n_8), .CO(n_9), .S(p_2[25]));
   FA_X1 i_10 (.A(p_0[26]), .B(p_1[26]), .CI(n_9), .CO(n_10), .S(p_2[26]));
   FA_X1 i_11 (.A(p_0[27]), .B(p_1[27]), .CI(n_10), .CO(n_11), .S(p_2[27]));
   FA_X1 i_12 (.A(p_0[28]), .B(p_1[28]), .CI(n_11), .CO(n_12), .S(p_2[28]));
   FA_X1 i_13 (.A(p_0[29]), .B(p_1[29]), .CI(n_12), .CO(n_13), .S(p_2[29]));
   FA_X1 i_14 (.A(p_0[30]), .B(p_1[30]), .CI(n_13), .CO(n_14), .S(p_2[30]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[31]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[31]), .B1(p_0[31]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[32]), .B(n_15), .Z(p_2[32]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[31]), .A3(n_16), .B1(p_0[31]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[31]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[31]), .ZN(n_18));
endmodule

module datapath__0_43(p_0, p_1, p_2);
   input [32:0]p_0;
   input [32:0]p_1;
   output [32:0]p_2;

   HA_X1 i_1 (.A(p_0[17]), .B(p_1[17]), .CO(n_1), .S(p_2[17]));
   FA_X1 i_2 (.A(p_0[18]), .B(p_1[18]), .CI(n_1), .CO(n_2), .S(p_2[18]));
   FA_X1 i_3 (.A(p_0[19]), .B(p_1[19]), .CI(n_2), .CO(n_3), .S(p_2[19]));
   FA_X1 i_4 (.A(p_0[20]), .B(p_1[20]), .CI(n_3), .CO(n_4), .S(p_2[20]));
   FA_X1 i_5 (.A(p_0[21]), .B(p_1[21]), .CI(n_4), .CO(n_5), .S(p_2[21]));
   FA_X1 i_6 (.A(p_0[22]), .B(p_1[22]), .CI(n_5), .CO(n_6), .S(p_2[22]));
   FA_X1 i_7 (.A(p_0[23]), .B(p_1[23]), .CI(n_6), .CO(n_7), .S(p_2[23]));
   FA_X1 i_8 (.A(p_0[24]), .B(p_1[24]), .CI(n_7), .CO(n_8), .S(p_2[24]));
   FA_X1 i_9 (.A(p_0[25]), .B(p_1[25]), .CI(n_8), .CO(n_9), .S(p_2[25]));
   FA_X1 i_10 (.A(p_0[26]), .B(p_1[26]), .CI(n_9), .CO(n_10), .S(p_2[26]));
   FA_X1 i_11 (.A(p_0[27]), .B(p_1[27]), .CI(n_10), .CO(n_11), .S(p_2[27]));
   FA_X1 i_12 (.A(p_0[28]), .B(p_1[28]), .CI(n_11), .CO(n_12), .S(p_2[28]));
   FA_X1 i_13 (.A(p_0[29]), .B(p_1[29]), .CI(n_12), .CO(n_13), .S(p_2[29]));
   FA_X1 i_14 (.A(p_0[30]), .B(p_1[30]), .CI(n_13), .CO(n_14), .S(p_2[30]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[31]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[31]), .B1(p_0[31]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[32]), .B(n_15), .Z(p_2[32]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[31]), .A3(n_16), .B1(p_0[31]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[31]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[31]), .ZN(n_18));
endmodule

module datapath__0_46(p_0, p_1, p_2);
   input [32:0]p_0;
   input [32:0]p_1;
   output [32:0]p_2;

   HA_X1 i_1 (.A(p_0[17]), .B(p_1[17]), .CO(n_1), .S(p_2[17]));
   FA_X1 i_2 (.A(p_0[18]), .B(p_1[18]), .CI(n_1), .CO(n_2), .S(p_2[18]));
   FA_X1 i_3 (.A(p_0[19]), .B(p_1[19]), .CI(n_2), .CO(n_3), .S(p_2[19]));
   FA_X1 i_4 (.A(p_0[20]), .B(p_1[20]), .CI(n_3), .CO(n_4), .S(p_2[20]));
   FA_X1 i_5 (.A(p_0[21]), .B(p_1[21]), .CI(n_4), .CO(n_5), .S(p_2[21]));
   FA_X1 i_6 (.A(p_0[22]), .B(p_1[22]), .CI(n_5), .CO(n_6), .S(p_2[22]));
   FA_X1 i_7 (.A(p_0[23]), .B(p_1[23]), .CI(n_6), .CO(n_7), .S(p_2[23]));
   FA_X1 i_8 (.A(p_0[24]), .B(p_1[24]), .CI(n_7), .CO(n_8), .S(p_2[24]));
   FA_X1 i_9 (.A(p_0[25]), .B(p_1[25]), .CI(n_8), .CO(n_9), .S(p_2[25]));
   FA_X1 i_10 (.A(p_0[26]), .B(p_1[26]), .CI(n_9), .CO(n_10), .S(p_2[26]));
   FA_X1 i_11 (.A(p_0[27]), .B(p_1[27]), .CI(n_10), .CO(n_11), .S(p_2[27]));
   FA_X1 i_12 (.A(p_0[28]), .B(p_1[28]), .CI(n_11), .CO(n_12), .S(p_2[28]));
   FA_X1 i_13 (.A(p_0[29]), .B(p_1[29]), .CI(n_12), .CO(n_13), .S(p_2[29]));
   FA_X1 i_14 (.A(p_0[30]), .B(p_1[30]), .CI(n_13), .CO(n_14), .S(p_2[30]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[31]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[31]), .B1(p_0[31]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[32]), .B(n_15), .Z(p_2[32]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[31]), .A3(n_16), .B1(p_0[31]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[31]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[31]), .ZN(n_18));
endmodule

module datapath__0_47(p_0, p_1, p_2);
   input [32:0]p_0;
   input [32:0]p_1;
   output [32:0]p_2;

   HA_X1 i_1 (.A(p_0[17]), .B(p_1[17]), .CO(n_1), .S(p_2[17]));
   FA_X1 i_2 (.A(p_0[18]), .B(p_1[18]), .CI(n_1), .CO(n_2), .S(p_2[18]));
   FA_X1 i_3 (.A(p_0[19]), .B(p_1[19]), .CI(n_2), .CO(n_3), .S(p_2[19]));
   FA_X1 i_4 (.A(p_0[20]), .B(p_1[20]), .CI(n_3), .CO(n_4), .S(p_2[20]));
   FA_X1 i_5 (.A(p_0[21]), .B(p_1[21]), .CI(n_4), .CO(n_5), .S(p_2[21]));
   FA_X1 i_6 (.A(p_0[22]), .B(p_1[22]), .CI(n_5), .CO(n_6), .S(p_2[22]));
   FA_X1 i_7 (.A(p_0[23]), .B(p_1[23]), .CI(n_6), .CO(n_7), .S(p_2[23]));
   FA_X1 i_8 (.A(p_0[24]), .B(p_1[24]), .CI(n_7), .CO(n_8), .S(p_2[24]));
   FA_X1 i_9 (.A(p_0[25]), .B(p_1[25]), .CI(n_8), .CO(n_9), .S(p_2[25]));
   FA_X1 i_10 (.A(p_0[26]), .B(p_1[26]), .CI(n_9), .CO(n_10), .S(p_2[26]));
   FA_X1 i_11 (.A(p_0[27]), .B(p_1[27]), .CI(n_10), .CO(n_11), .S(p_2[27]));
   FA_X1 i_12 (.A(p_0[28]), .B(p_1[28]), .CI(n_11), .CO(n_12), .S(p_2[28]));
   FA_X1 i_13 (.A(p_0[29]), .B(p_1[29]), .CI(n_12), .CO(n_13), .S(p_2[29]));
   FA_X1 i_14 (.A(p_0[30]), .B(p_1[30]), .CI(n_13), .CO(n_14), .S(p_2[30]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[31]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[31]), .B1(p_0[31]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[32]), .B(n_15), .Z(p_2[32]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[31]), .A3(n_16), .B1(p_0[31]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[31]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[31]), .ZN(n_18));
endmodule

module datapath__0_50(p_0, p_1, p_2);
   input [32:0]p_0;
   input [32:0]p_1;
   output [32:0]p_2;

   HA_X1 i_1 (.A(p_0[17]), .B(p_1[17]), .CO(n_1), .S(p_2[17]));
   FA_X1 i_2 (.A(p_0[18]), .B(p_1[18]), .CI(n_1), .CO(n_2), .S(p_2[18]));
   FA_X1 i_3 (.A(p_0[19]), .B(p_1[19]), .CI(n_2), .CO(n_3), .S(p_2[19]));
   FA_X1 i_4 (.A(p_0[20]), .B(p_1[20]), .CI(n_3), .CO(n_4), .S(p_2[20]));
   FA_X1 i_5 (.A(p_0[21]), .B(p_1[21]), .CI(n_4), .CO(n_5), .S(p_2[21]));
   FA_X1 i_6 (.A(p_0[22]), .B(p_1[22]), .CI(n_5), .CO(n_6), .S(p_2[22]));
   FA_X1 i_7 (.A(p_0[23]), .B(p_1[23]), .CI(n_6), .CO(n_7), .S(p_2[23]));
   FA_X1 i_8 (.A(p_0[24]), .B(p_1[24]), .CI(n_7), .CO(n_8), .S(p_2[24]));
   FA_X1 i_9 (.A(p_0[25]), .B(p_1[25]), .CI(n_8), .CO(n_9), .S(p_2[25]));
   FA_X1 i_10 (.A(p_0[26]), .B(p_1[26]), .CI(n_9), .CO(n_10), .S(p_2[26]));
   FA_X1 i_11 (.A(p_0[27]), .B(p_1[27]), .CI(n_10), .CO(n_11), .S(p_2[27]));
   FA_X1 i_12 (.A(p_0[28]), .B(p_1[28]), .CI(n_11), .CO(n_12), .S(p_2[28]));
   FA_X1 i_13 (.A(p_0[29]), .B(p_1[29]), .CI(n_12), .CO(n_13), .S(p_2[29]));
   FA_X1 i_14 (.A(p_0[30]), .B(p_1[30]), .CI(n_13), .CO(n_14), .S(p_2[30]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[31]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[31]), .B1(p_0[31]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[32]), .B(n_15), .Z(p_2[32]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[31]), .A3(n_16), .B1(p_0[31]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[31]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[31]), .ZN(n_18));
endmodule

module datapath__0_51(p_0, p_1, p_2);
   input [32:0]p_0;
   input [32:0]p_1;
   output [32:0]p_2;

   HA_X1 i_1 (.A(p_0[17]), .B(p_1[17]), .CO(n_1), .S(p_2[17]));
   FA_X1 i_2 (.A(p_0[18]), .B(p_1[18]), .CI(n_1), .CO(n_2), .S(p_2[18]));
   FA_X1 i_3 (.A(p_0[19]), .B(p_1[19]), .CI(n_2), .CO(n_3), .S(p_2[19]));
   FA_X1 i_4 (.A(p_0[20]), .B(p_1[20]), .CI(n_3), .CO(n_4), .S(p_2[20]));
   FA_X1 i_5 (.A(p_0[21]), .B(p_1[21]), .CI(n_4), .CO(n_5), .S(p_2[21]));
   FA_X1 i_6 (.A(p_0[22]), .B(p_1[22]), .CI(n_5), .CO(n_6), .S(p_2[22]));
   FA_X1 i_7 (.A(p_0[23]), .B(p_1[23]), .CI(n_6), .CO(n_7), .S(p_2[23]));
   FA_X1 i_8 (.A(p_0[24]), .B(p_1[24]), .CI(n_7), .CO(n_8), .S(p_2[24]));
   FA_X1 i_9 (.A(p_0[25]), .B(p_1[25]), .CI(n_8), .CO(n_9), .S(p_2[25]));
   FA_X1 i_10 (.A(p_0[26]), .B(p_1[26]), .CI(n_9), .CO(n_10), .S(p_2[26]));
   FA_X1 i_11 (.A(p_0[27]), .B(p_1[27]), .CI(n_10), .CO(n_11), .S(p_2[27]));
   FA_X1 i_12 (.A(p_0[28]), .B(p_1[28]), .CI(n_11), .CO(n_12), .S(p_2[28]));
   FA_X1 i_13 (.A(p_0[29]), .B(p_1[29]), .CI(n_12), .CO(n_13), .S(p_2[29]));
   FA_X1 i_14 (.A(p_0[30]), .B(p_1[30]), .CI(n_13), .CO(n_14), .S(p_2[30]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[31]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[31]), .B1(p_0[31]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[32]), .B(n_15), .Z(p_2[32]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[31]), .A3(n_16), .B1(p_0[31]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[31]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[31]), .ZN(n_18));
endmodule

module datapath__0_54(p_0, p_1, p_2);
   input [32:0]p_0;
   input [32:0]p_1;
   output [32:0]p_2;

   HA_X1 i_1 (.A(p_0[17]), .B(p_1[17]), .CO(n_1), .S(p_2[17]));
   FA_X1 i_2 (.A(p_0[18]), .B(p_1[18]), .CI(n_1), .CO(n_2), .S(p_2[18]));
   FA_X1 i_3 (.A(p_0[19]), .B(p_1[19]), .CI(n_2), .CO(n_3), .S(p_2[19]));
   FA_X1 i_4 (.A(p_0[20]), .B(p_1[20]), .CI(n_3), .CO(n_4), .S(p_2[20]));
   FA_X1 i_5 (.A(p_0[21]), .B(p_1[21]), .CI(n_4), .CO(n_5), .S(p_2[21]));
   FA_X1 i_6 (.A(p_0[22]), .B(p_1[22]), .CI(n_5), .CO(n_6), .S(p_2[22]));
   FA_X1 i_7 (.A(p_0[23]), .B(p_1[23]), .CI(n_6), .CO(n_7), .S(p_2[23]));
   FA_X1 i_8 (.A(p_0[24]), .B(p_1[24]), .CI(n_7), .CO(n_8), .S(p_2[24]));
   FA_X1 i_9 (.A(p_0[25]), .B(p_1[25]), .CI(n_8), .CO(n_9), .S(p_2[25]));
   FA_X1 i_10 (.A(p_0[26]), .B(p_1[26]), .CI(n_9), .CO(n_10), .S(p_2[26]));
   FA_X1 i_11 (.A(p_0[27]), .B(p_1[27]), .CI(n_10), .CO(n_11), .S(p_2[27]));
   FA_X1 i_12 (.A(p_0[28]), .B(p_1[28]), .CI(n_11), .CO(n_12), .S(p_2[28]));
   FA_X1 i_13 (.A(p_0[29]), .B(p_1[29]), .CI(n_12), .CO(n_13), .S(p_2[29]));
   FA_X1 i_14 (.A(p_0[30]), .B(p_1[30]), .CI(n_13), .CO(n_14), .S(p_2[30]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[31]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[31]), .B1(p_0[31]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[32]), .B(n_15), .Z(p_2[32]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[31]), .A3(n_16), .B1(p_0[31]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[31]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[31]), .ZN(n_18));
endmodule

module datapath__0_55(p_0, p_1, p_2);
   input [32:0]p_0;
   input [32:0]p_1;
   output [32:0]p_2;

   HA_X1 i_1 (.A(p_0[17]), .B(p_1[17]), .CO(n_1), .S(p_2[17]));
   FA_X1 i_2 (.A(p_0[18]), .B(p_1[18]), .CI(n_1), .CO(n_2), .S(p_2[18]));
   FA_X1 i_3 (.A(p_0[19]), .B(p_1[19]), .CI(n_2), .CO(n_3), .S(p_2[19]));
   FA_X1 i_4 (.A(p_0[20]), .B(p_1[20]), .CI(n_3), .CO(n_4), .S(p_2[20]));
   FA_X1 i_5 (.A(p_0[21]), .B(p_1[21]), .CI(n_4), .CO(n_5), .S(p_2[21]));
   FA_X1 i_6 (.A(p_0[22]), .B(p_1[22]), .CI(n_5), .CO(n_6), .S(p_2[22]));
   FA_X1 i_7 (.A(p_0[23]), .B(p_1[23]), .CI(n_6), .CO(n_7), .S(p_2[23]));
   FA_X1 i_8 (.A(p_0[24]), .B(p_1[24]), .CI(n_7), .CO(n_8), .S(p_2[24]));
   FA_X1 i_9 (.A(p_0[25]), .B(p_1[25]), .CI(n_8), .CO(n_9), .S(p_2[25]));
   FA_X1 i_10 (.A(p_0[26]), .B(p_1[26]), .CI(n_9), .CO(n_10), .S(p_2[26]));
   FA_X1 i_11 (.A(p_0[27]), .B(p_1[27]), .CI(n_10), .CO(n_11), .S(p_2[27]));
   FA_X1 i_12 (.A(p_0[28]), .B(p_1[28]), .CI(n_11), .CO(n_12), .S(p_2[28]));
   FA_X1 i_13 (.A(p_0[29]), .B(p_1[29]), .CI(n_12), .CO(n_13), .S(p_2[29]));
   FA_X1 i_14 (.A(p_0[30]), .B(p_1[30]), .CI(n_13), .CO(n_14), .S(p_2[30]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[31]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[31]), .B1(p_0[31]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[32]), .B(n_15), .Z(p_2[32]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[31]), .A3(n_16), .B1(p_0[31]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[31]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[31]), .ZN(n_18));
endmodule

module datapath__0_58(p_0, p_1, p_2);
   input [32:0]p_0;
   input [32:0]p_1;
   output [32:0]p_2;

   HA_X1 i_1 (.A(p_0[17]), .B(p_1[17]), .CO(n_1), .S(p_2[17]));
   FA_X1 i_2 (.A(p_0[18]), .B(p_1[18]), .CI(n_1), .CO(n_2), .S(p_2[18]));
   FA_X1 i_3 (.A(p_0[19]), .B(p_1[19]), .CI(n_2), .CO(n_3), .S(p_2[19]));
   FA_X1 i_4 (.A(p_0[20]), .B(p_1[20]), .CI(n_3), .CO(n_4), .S(p_2[20]));
   FA_X1 i_5 (.A(p_0[21]), .B(p_1[21]), .CI(n_4), .CO(n_5), .S(p_2[21]));
   FA_X1 i_6 (.A(p_0[22]), .B(p_1[22]), .CI(n_5), .CO(n_6), .S(p_2[22]));
   FA_X1 i_7 (.A(p_0[23]), .B(p_1[23]), .CI(n_6), .CO(n_7), .S(p_2[23]));
   FA_X1 i_8 (.A(p_0[24]), .B(p_1[24]), .CI(n_7), .CO(n_8), .S(p_2[24]));
   FA_X1 i_9 (.A(p_0[25]), .B(p_1[25]), .CI(n_8), .CO(n_9), .S(p_2[25]));
   FA_X1 i_10 (.A(p_0[26]), .B(p_1[26]), .CI(n_9), .CO(n_10), .S(p_2[26]));
   FA_X1 i_11 (.A(p_0[27]), .B(p_1[27]), .CI(n_10), .CO(n_11), .S(p_2[27]));
   FA_X1 i_12 (.A(p_0[28]), .B(p_1[28]), .CI(n_11), .CO(n_12), .S(p_2[28]));
   FA_X1 i_13 (.A(p_0[29]), .B(p_1[29]), .CI(n_12), .CO(n_13), .S(p_2[29]));
   FA_X1 i_14 (.A(p_0[30]), .B(p_1[30]), .CI(n_13), .CO(n_14), .S(p_2[30]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[31]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[31]), .B1(p_0[31]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[32]), .B(n_15), .Z(p_2[32]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[31]), .A3(n_16), .B1(p_0[31]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[31]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[31]), .ZN(n_18));
endmodule

module datapath__0_59(p_0, p_1, p_2);
   input [32:0]p_0;
   input [32:0]p_1;
   output [32:0]p_2;

   HA_X1 i_1 (.A(p_0[17]), .B(p_1[17]), .CO(n_1), .S(p_2[17]));
   FA_X1 i_2 (.A(p_0[18]), .B(p_1[18]), .CI(n_1), .CO(n_2), .S(p_2[18]));
   FA_X1 i_3 (.A(p_0[19]), .B(p_1[19]), .CI(n_2), .CO(n_3), .S(p_2[19]));
   FA_X1 i_4 (.A(p_0[20]), .B(p_1[20]), .CI(n_3), .CO(n_4), .S(p_2[20]));
   FA_X1 i_5 (.A(p_0[21]), .B(p_1[21]), .CI(n_4), .CO(n_5), .S(p_2[21]));
   FA_X1 i_6 (.A(p_0[22]), .B(p_1[22]), .CI(n_5), .CO(n_6), .S(p_2[22]));
   FA_X1 i_7 (.A(p_0[23]), .B(p_1[23]), .CI(n_6), .CO(n_7), .S(p_2[23]));
   FA_X1 i_8 (.A(p_0[24]), .B(p_1[24]), .CI(n_7), .CO(n_8), .S(p_2[24]));
   FA_X1 i_9 (.A(p_0[25]), .B(p_1[25]), .CI(n_8), .CO(n_9), .S(p_2[25]));
   FA_X1 i_10 (.A(p_0[26]), .B(p_1[26]), .CI(n_9), .CO(n_10), .S(p_2[26]));
   FA_X1 i_11 (.A(p_0[27]), .B(p_1[27]), .CI(n_10), .CO(n_11), .S(p_2[27]));
   FA_X1 i_12 (.A(p_0[28]), .B(p_1[28]), .CI(n_11), .CO(n_12), .S(p_2[28]));
   FA_X1 i_13 (.A(p_0[29]), .B(p_1[29]), .CI(n_12), .CO(n_13), .S(p_2[29]));
   FA_X1 i_14 (.A(p_0[30]), .B(p_1[30]), .CI(n_13), .CO(n_14), .S(p_2[30]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_2[31]));
   OAI22_X1 i_15 (.A1(n_18), .A2(p_1[31]), .B1(p_0[31]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(p_0[32]), .B(n_15), .Z(p_2[32]));
   OAI33_X1 i_17 (.A1(n_18), .A2(p_1[31]), .A3(n_16), .B1(p_0[31]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(p_1[31]), .ZN(n_17));
   INV_X1 i_20 (.A(p_0[31]), .ZN(n_18));
endmodule

module Booth_Multiplier(multiplicand, multiplier, product);
   input [15:0]multiplicand;
   input [15:0]multiplier;
   output [31:0]product;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_215;
   wire n_0_216;
   wire n_0_217;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_230;
   wire n_0_231;
   wire n_0_232;
   wire n_0_233;
   wire n_0_234;
   wire n_0_235;
   wire n_0_236;
   wire n_0_237;
   wire n_0_238;
   wire n_0_239;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_248;
   wire n_0_249;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_256;
   wire n_0_257;
   wire n_0_258;
   wire n_0_259;
   wire n_0_260;
   wire n_0_261;
   wire n_0_262;
   wire n_0_263;
   wire n_0_264;
   wire n_0_265;
   wire n_0_266;
   wire n_0_267;
   wire n_0_268;
   wire n_0_269;
   wire n_0_270;
   wire n_0_271;
   wire n_0_272;
   wire n_0_273;
   wire n_0_274;
   wire n_0_275;
   wire n_0_276;
   wire n_0_277;
   wire n_0_278;
   wire n_0_279;
   wire n_0_280;
   wire n_0_281;
   wire n_0_282;
   wire n_0_283;
   wire n_0_284;
   wire n_0_285;
   wire n_0_286;
   wire n_0_287;
   wire n_0_288;
   wire n_0_289;
   wire n_0_290;
   wire n_0_291;
   wire n_0_292;
   wire n_0_293;
   wire n_0_294;
   wire n_0_295;
   wire n_0_296;
   wire n_0_297;
   wire n_0_298;
   wire n_0_299;
   wire n_0_300;
   wire n_0_301;
   wire n_0_302;
   wire n_0_303;
   wire n_0_304;
   wire n_0_305;
   wire n_0_306;
   wire n_0_307;
   wire n_0_308;
   wire n_0_309;
   wire n_0_310;
   wire n_0_311;
   wire n_0_312;
   wire n_0_313;
   wire n_0_314;
   wire n_0_315;
   wire n_0_316;
   wire n_0_317;
   wire n_0_318;
   wire n_0_319;
   wire n_0_320;
   wire n_0_321;
   wire n_0_322;
   wire n_0_323;
   wire n_0_324;
   wire n_0_325;
   wire n_0_326;
   wire n_0_327;
   wire n_0_328;
   wire n_0_329;
   wire n_0_330;
   wire n_0_331;
   wire n_0_332;
   wire n_0_333;
   wire n_0_334;
   wire n_0_335;
   wire n_0_336;
   wire n_0_337;
   wire n_0_338;
   wire n_0_339;
   wire n_0_340;
   wire n_0_341;
   wire n_0_342;
   wire n_0_343;
   wire n_0_344;
   wire n_0_345;
   wire n_0_346;
   wire n_0_347;
   wire n_0_348;
   wire n_0_349;
   wire n_0_350;
   wire n_0_351;
   wire n_0_352;
   wire n_0_353;
   wire n_0_354;
   wire n_0_355;
   wire n_0_356;
   wire n_0_357;
   wire n_0_358;
   wire n_0_359;
   wire n_0_360;
   wire n_0_361;
   wire n_0_362;
   wire n_0_363;
   wire n_0_364;
   wire n_0_365;
   wire n_0_366;
   wire n_0_367;
   wire n_0_368;
   wire n_0_369;
   wire n_0_370;
   wire n_0_371;
   wire n_0_372;
   wire n_0_373;
   wire n_0_374;
   wire n_0_375;
   wire n_0_376;
   wire n_0_377;
   wire n_0_378;
   wire n_0_379;
   wire n_0_380;
   wire n_0_381;
   wire n_0_382;
   wire n_0_383;
   wire n_0_384;
   wire n_0_385;
   wire n_0_386;
   wire n_0_387;
   wire n_0_388;
   wire n_0_389;
   wire n_0_390;
   wire n_0_391;
   wire n_0_392;
   wire n_0_393;
   wire n_0_394;
   wire n_0_395;
   wire n_0_396;
   wire n_0_397;
   wire n_0_398;
   wire n_0_399;
   wire n_0_400;
   wire n_0_401;
   wire n_0_402;
   wire n_0_403;
   wire n_0_404;
   wire n_0_405;
   wire n_0_406;
   wire n_0_407;
   wire n_0_408;
   wire n_0_409;
   wire n_0_410;
   wire n_0_411;
   wire n_0_412;
   wire n_0_413;
   wire n_0_414;
   wire n_0_415;
   wire n_0_416;
   wire n_0_417;
   wire n_0_418;
   wire n_0_419;
   wire n_0_420;
   wire n_0_421;
   wire n_0_422;
   wire n_0_423;
   wire n_0_424;
   wire n_0_425;
   wire n_0_426;
   wire n_0_427;
   wire n_0_428;
   wire n_0_429;
   wire n_0_430;
   wire n_0_431;
   wire n_0_432;
   wire n_0_433;
   wire n_0_434;
   wire n_0_435;
   wire n_0_436;
   wire n_0_437;
   wire n_0_438;
   wire n_0_439;
   wire n_0_440;
   wire n_0_441;
   wire n_0_442;
   wire n_0_443;
   wire n_0_444;
   wire n_0_445;
   wire n_0_446;
   wire n_0_447;
   wire n_0_448;
   wire n_0_449;
   wire n_0_450;
   wire n_0_451;
   wire n_0_452;
   wire n_0_453;
   wire n_0_454;
   wire n_0_455;
   wire n_0_456;
   wire n_0_457;
   wire n_0_458;
   wire n_0_459;
   wire n_0_460;
   wire n_0_461;
   wire n_0_462;
   wire n_0_463;
   wire n_0_464;
   wire n_0_465;
   wire n_0_466;
   wire n_0_467;
   wire n_0_468;
   wire n_0_469;
   wire n_0_470;
   wire n_0_471;
   wire n_0_472;
   wire n_0_473;
   wire n_0_474;
   wire n_0_475;
   wire n_0_476;
   wire n_0_477;
   wire n_0_478;
   wire n_0_479;
   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_0_7;
   wire n_0_0_8;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_480;
   wire n_0_0_21;
   wire n_0_481;
   wire n_0_0_22;
   wire n_0_482;
   wire n_0_0_23;
   wire n_0_483;
   wire n_0_0_24;
   wire n_0_484;
   wire n_0_0_25;
   wire n_0_485;
   wire n_0_0_26;
   wire n_0_486;
   wire n_0_0_27;
   wire n_0_487;
   wire n_0_0_28;
   wire n_0_488;
   wire n_0_0_29;
   wire n_0_489;
   wire n_0_0_30;
   wire n_0_490;
   wire n_0_0_31;
   wire n_0_491;
   wire n_0_0_32;
   wire n_0_492;
   wire n_0_0_33;
   wire n_0_493;
   wire n_0_0_34;
   wire n_0_494;
   wire n_0_0_35;
   wire n_0_0_36;
   wire n_0_0_37;
   wire n_0_0_38;
   wire n_0_0_39;
   wire n_0_0_40;
   wire n_0_495;
   wire n_0_0_41;
   wire n_0_496;
   wire n_0_0_42;
   wire n_0_497;
   wire n_0_0_43;
   wire n_0_498;
   wire n_0_0_44;
   wire n_0_499;
   wire n_0_0_45;
   wire n_0_500;
   wire n_0_0_46;
   wire n_0_501;
   wire n_0_0_47;
   wire n_0_502;
   wire n_0_0_48;
   wire n_0_503;
   wire n_0_0_49;
   wire n_0_504;
   wire n_0_0_50;
   wire n_0_505;
   wire n_0_0_51;
   wire n_0_506;
   wire n_0_0_52;
   wire n_0_507;
   wire n_0_0_53;
   wire n_0_508;
   wire n_0_0_54;
   wire n_0_509;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_510;
   wire n_0_0_61;
   wire n_0_511;
   wire n_0_0_62;
   wire n_0_512;
   wire n_0_0_63;
   wire n_0_513;
   wire n_0_0_64;
   wire n_0_514;
   wire n_0_0_65;
   wire n_0_515;
   wire n_0_0_66;
   wire n_0_516;
   wire n_0_0_67;
   wire n_0_517;
   wire n_0_0_68;
   wire n_0_518;
   wire n_0_0_69;
   wire n_0_519;
   wire n_0_0_70;
   wire n_0_520;
   wire n_0_0_71;
   wire n_0_521;
   wire n_0_0_72;
   wire n_0_522;
   wire n_0_0_73;
   wire n_0_523;
   wire n_0_0_74;
   wire n_0_524;
   wire n_0_0_75;
   wire n_0_0_76;
   wire n_0_0_77;
   wire n_0_0_78;
   wire n_0_0_79;
   wire n_0_0_80;
   wire n_0_525;
   wire n_0_0_81;
   wire n_0_526;
   wire n_0_0_82;
   wire n_0_527;
   wire n_0_0_83;
   wire n_0_528;
   wire n_0_0_84;
   wire n_0_529;
   wire n_0_0_85;
   wire n_0_530;
   wire n_0_0_86;
   wire n_0_531;
   wire n_0_0_87;
   wire n_0_532;
   wire n_0_0_88;
   wire n_0_533;
   wire n_0_0_89;
   wire n_0_534;
   wire n_0_0_90;
   wire n_0_535;
   wire n_0_0_91;
   wire n_0_536;
   wire n_0_0_92;
   wire n_0_537;
   wire n_0_0_93;
   wire n_0_538;
   wire n_0_0_94;
   wire n_0_539;
   wire n_0_0_95;
   wire n_0_0_96;
   wire n_0_0_97;
   wire n_0_0_98;
   wire n_0_0_99;
   wire n_0_0_100;
   wire n_0_540;
   wire n_0_0_101;
   wire n_0_541;
   wire n_0_0_102;
   wire n_0_542;
   wire n_0_0_103;
   wire n_0_543;
   wire n_0_0_104;
   wire n_0_544;
   wire n_0_0_105;
   wire n_0_545;
   wire n_0_0_106;
   wire n_0_546;
   wire n_0_0_107;
   wire n_0_547;
   wire n_0_0_108;
   wire n_0_548;
   wire n_0_0_109;
   wire n_0_549;
   wire n_0_0_110;
   wire n_0_550;
   wire n_0_0_111;
   wire n_0_551;
   wire n_0_0_112;
   wire n_0_552;
   wire n_0_0_113;
   wire n_0_553;
   wire n_0_0_114;
   wire n_0_554;
   wire n_0_0_115;
   wire n_0_0_116;
   wire n_0_0_117;
   wire n_0_0_118;
   wire n_0_0_119;
   wire n_0_0_120;
   wire n_0_555;
   wire n_0_0_121;
   wire n_0_556;
   wire n_0_0_122;
   wire n_0_557;
   wire n_0_0_123;
   wire n_0_558;
   wire n_0_0_124;
   wire n_0_559;
   wire n_0_0_125;
   wire n_0_560;
   wire n_0_0_126;
   wire n_0_561;
   wire n_0_0_127;
   wire n_0_562;
   wire n_0_0_128;
   wire n_0_563;
   wire n_0_0_129;
   wire n_0_564;
   wire n_0_0_130;
   wire n_0_565;
   wire n_0_0_131;
   wire n_0_566;
   wire n_0_0_132;
   wire n_0_567;
   wire n_0_0_133;
   wire n_0_568;
   wire n_0_0_134;
   wire n_0_569;
   wire n_0_0_135;
   wire n_0_0_136;
   wire n_0_0_137;
   wire n_0_0_138;
   wire n_0_0_139;
   wire n_0_0_140;
   wire n_0_570;
   wire n_0_0_141;
   wire n_0_571;
   wire n_0_0_142;
   wire n_0_572;
   wire n_0_0_143;
   wire n_0_573;
   wire n_0_0_144;
   wire n_0_574;
   wire n_0_0_145;
   wire n_0_575;
   wire n_0_0_146;
   wire n_0_576;
   wire n_0_0_147;
   wire n_0_577;
   wire n_0_0_148;
   wire n_0_578;
   wire n_0_0_149;
   wire n_0_579;
   wire n_0_0_150;
   wire n_0_580;
   wire n_0_0_151;
   wire n_0_581;
   wire n_0_0_152;
   wire n_0_582;
   wire n_0_0_153;
   wire n_0_583;
   wire n_0_0_154;
   wire n_0_584;
   wire n_0_0_155;
   wire n_0_0_156;
   wire n_0_0_157;
   wire n_0_0_158;
   wire n_0_0_159;
   wire n_0_0_160;
   wire n_0_585;
   wire n_0_0_161;
   wire n_0_586;
   wire n_0_0_162;
   wire n_0_587;
   wire n_0_0_163;
   wire n_0_588;
   wire n_0_0_164;
   wire n_0_589;
   wire n_0_0_165;
   wire n_0_590;
   wire n_0_0_166;
   wire n_0_591;
   wire n_0_0_167;
   wire n_0_592;
   wire n_0_0_168;
   wire n_0_593;
   wire n_0_0_169;
   wire n_0_594;
   wire n_0_0_170;
   wire n_0_595;
   wire n_0_0_171;
   wire n_0_596;
   wire n_0_0_172;
   wire n_0_597;
   wire n_0_0_173;
   wire n_0_598;
   wire n_0_0_174;
   wire n_0_599;
   wire n_0_0_175;
   wire n_0_0_176;
   wire n_0_0_177;
   wire n_0_0_178;
   wire n_0_0_179;
   wire n_0_0_180;
   wire n_0_600;
   wire n_0_0_181;
   wire n_0_601;
   wire n_0_0_182;
   wire n_0_602;
   wire n_0_0_183;
   wire n_0_603;
   wire n_0_0_184;
   wire n_0_604;
   wire n_0_0_185;
   wire n_0_605;
   wire n_0_0_186;
   wire n_0_606;
   wire n_0_0_187;
   wire n_0_607;
   wire n_0_0_188;
   wire n_0_608;
   wire n_0_0_189;
   wire n_0_609;
   wire n_0_0_190;
   wire n_0_610;
   wire n_0_0_191;
   wire n_0_611;
   wire n_0_0_192;
   wire n_0_612;
   wire n_0_0_193;
   wire n_0_613;
   wire n_0_0_194;
   wire n_0_614;
   wire n_0_0_195;
   wire n_0_0_196;
   wire n_0_0_197;
   wire n_0_0_198;
   wire n_0_0_199;
   wire n_0_0_200;
   wire n_0_615;
   wire n_0_0_201;
   wire n_0_616;
   wire n_0_0_202;
   wire n_0_617;
   wire n_0_0_203;
   wire n_0_618;
   wire n_0_0_204;
   wire n_0_619;
   wire n_0_0_205;
   wire n_0_620;
   wire n_0_0_206;
   wire n_0_621;
   wire n_0_0_207;
   wire n_0_622;
   wire n_0_0_208;
   wire n_0_623;
   wire n_0_0_209;
   wire n_0_624;
   wire n_0_0_210;
   wire n_0_625;
   wire n_0_0_211;
   wire n_0_626;
   wire n_0_0_212;
   wire n_0_627;
   wire n_0_0_213;
   wire n_0_628;
   wire n_0_0_214;
   wire n_0_629;
   wire n_0_0_215;
   wire n_0_0_216;
   wire n_0_0_217;
   wire n_0_0_218;
   wire n_0_0_219;
   wire n_0_0_220;
   wire n_0_630;
   wire n_0_0_221;
   wire n_0_631;
   wire n_0_0_222;
   wire n_0_632;
   wire n_0_0_223;
   wire n_0_633;
   wire n_0_0_224;
   wire n_0_634;
   wire n_0_0_225;
   wire n_0_635;
   wire n_0_0_226;
   wire n_0_636;
   wire n_0_0_227;
   wire n_0_637;
   wire n_0_0_228;
   wire n_0_638;
   wire n_0_0_229;
   wire n_0_639;
   wire n_0_0_230;
   wire n_0_640;
   wire n_0_0_231;
   wire n_0_641;
   wire n_0_0_232;
   wire n_0_642;
   wire n_0_0_233;
   wire n_0_643;
   wire n_0_0_234;
   wire n_0_644;
   wire n_0_0_235;
   wire n_0_0_236;
   wire n_0_0_237;
   wire n_0_0_238;
   wire n_0_0_239;
   wire n_0_0_240;
   wire n_0_645;
   wire n_0_0_241;
   wire n_0_646;
   wire n_0_0_242;
   wire n_0_647;
   wire n_0_0_243;
   wire n_0_648;
   wire n_0_0_244;
   wire n_0_649;
   wire n_0_0_245;
   wire n_0_650;
   wire n_0_0_246;
   wire n_0_651;
   wire n_0_0_247;
   wire n_0_652;
   wire n_0_0_248;
   wire n_0_653;
   wire n_0_0_249;
   wire n_0_654;
   wire n_0_0_250;
   wire n_0_655;
   wire n_0_0_251;
   wire n_0_656;
   wire n_0_0_252;
   wire n_0_657;
   wire n_0_0_253;
   wire n_0_658;
   wire n_0_0_254;
   wire n_0_659;
   wire n_0_0_255;
   wire n_0_0_256;
   wire n_0_0_257;
   wire n_0_0_258;
   wire n_0_0_259;
   wire n_0_0_260;
   wire n_0_660;
   wire n_0_0_261;
   wire n_0_661;
   wire n_0_0_262;
   wire n_0_662;
   wire n_0_0_263;
   wire n_0_663;
   wire n_0_0_264;
   wire n_0_664;
   wire n_0_0_265;
   wire n_0_665;
   wire n_0_0_266;
   wire n_0_666;
   wire n_0_0_267;
   wire n_0_667;
   wire n_0_0_268;
   wire n_0_668;
   wire n_0_0_269;
   wire n_0_669;
   wire n_0_0_270;
   wire n_0_670;
   wire n_0_0_271;
   wire n_0_671;
   wire n_0_0_272;
   wire n_0_672;
   wire n_0_0_273;
   wire n_0_673;
   wire n_0_0_274;
   wire n_0_674;
   wire n_0_0_275;
   wire n_0_0_276;
   wire n_0_0_277;
   wire n_0_0_278;
   wire n_0_0_279;
   wire n_0_0_280;
   wire n_0_675;
   wire n_0_0_281;
   wire n_0_676;
   wire n_0_0_282;
   wire n_0_677;
   wire n_0_0_283;
   wire n_0_678;
   wire n_0_0_284;
   wire n_0_679;
   wire n_0_0_285;
   wire n_0_680;
   wire n_0_0_286;
   wire n_0_681;
   wire n_0_0_287;
   wire n_0_682;
   wire n_0_0_288;
   wire n_0_683;
   wire n_0_0_289;
   wire n_0_684;
   wire n_0_0_290;
   wire n_0_685;
   wire n_0_0_291;
   wire n_0_686;
   wire n_0_0_292;
   wire n_0_687;
   wire n_0_0_293;
   wire n_0_688;
   wire n_0_0_294;
   wire n_0_689;
   wire n_0_0_295;
   wire n_0_0_296;
   wire n_0_0_297;
   wire n_0_0_298;
   wire n_0_0_299;
   wire n_0_690;
   wire n_0_691;
   wire n_0_692;
   wire n_0_693;
   wire n_0_694;
   wire n_0_695;
   wire n_0_696;
   wire n_0_697;
   wire n_0_698;
   wire n_0_699;
   wire n_0_700;
   wire n_0_701;
   wire n_0_702;
   wire n_0_703;
   wire n_0_704;
   wire n_0_705;
   wire n_0_706;
   wire n_0_707;
   wire n_0_708;
   wire n_0_709;
   wire n_0_710;
   wire n_0_711;
   wire n_0_712;
   wire n_0_713;
   wire n_0_714;
   wire n_0_715;
   wire n_0_716;
   wire n_0_717;
   wire n_0_718;
   wire n_0_719;
   wire n_0_0_300;
   wire n_0_0_301;
   wire n_0_0_302;
   wire n_0_0_303;
   wire n_0_0_304;
   wire n_0_0_305;
   wire n_0_0_306;
   wire n_0_0_307;
   wire n_0_0_308;
   wire n_0_0_309;
   wire n_0_0_310;
   wire n_0_0_311;
   wire n_0_0_312;
   wire n_0_0_313;
   wire n_0_0_314;
   wire n_0_0_315;
   wire n_0_0_316;
   wire n_0_0_317;
   wire n_0_0_318;
   wire n_0_0_319;
   wire n_0_0_320;
   wire n_0_0_321;
   wire n_0_0_322;
   wire n_0_0_323;
   wire n_0_0_324;
   wire n_0_0_325;
   wire n_0_0_326;
   wire n_0_0_327;
   wire n_0_0_328;
   wire n_0_0_329;
   wire n_0_0_330;
   wire n_0_0_331;
   wire n_0_0_332;
   wire n_0_0_333;
   wire n_0_0_334;
   wire n_0_0_335;
   wire n_0_0_336;
   wire n_0_0_337;
   wire n_0_0_338;
   wire n_0_0_339;
   wire n_0_0_340;
   wire n_0_0_341;

   assign product[31] = product[30];

   datapath__0_2 i_0_2 (.p_0({n_0_719, n_0_718, n_0_717, n_0_716, n_0_715, 
      n_0_714, n_0_713, n_0_712, n_0_711, n_0_710, n_0_709, n_0_708, n_0_707, 
      n_0_706, n_0_705, multiplicand[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
      .p_1({uc_0, n_0_704, n_0_703, n_0_702, n_0_701, n_0_700, n_0_699, n_0_698, 
      n_0_697, n_0_696, n_0_695, n_0_694, n_0_693, n_0_692, n_0_691, n_0_690, 
      uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, uc_7, uc_8, uc_9, uc_10, uc_11, uc_12, 
      uc_13, uc_14, uc_15, uc_16, uc_17}), .p_2({n_0_15, n_0_14, n_0_13, n_0_12, 
      n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2, 
      n_0_1, n_0_0, uc_18, uc_19, uc_20, uc_21, uc_22, uc_23, uc_24, uc_25, 
      uc_26, uc_27, uc_28, uc_29, uc_30, uc_31, uc_32, uc_33, uc_34}));
   datapath__0_3 i_0_3 (.p_0({multiplicand[15], multiplicand[14], 
      multiplicand[13], multiplicand[12], multiplicand[11], multiplicand[10], 
      multiplicand[9], multiplicand[8], multiplicand[7], multiplicand[6], 
      multiplicand[5], multiplicand[4], multiplicand[3], multiplicand[2], 
      multiplicand[1], multiplicand[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .p_1({uc_35, 
      n_0_704, n_0_703, n_0_702, n_0_701, n_0_700, n_0_699, n_0_698, n_0_697, 
      n_0_696, n_0_695, n_0_694, n_0_693, n_0_692, n_0_691, n_0_690, uc_36, 
      uc_37, uc_38, uc_39, uc_40, uc_41, uc_42, uc_43, uc_44, uc_45, uc_46, 
      uc_47, uc_48, uc_49, uc_50, uc_51, uc_52}), .p_2({n_0_31, n_0_30, n_0_29, 
      n_0_28, n_0_27, n_0_26, n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, 
      n_0_19, n_0_18, n_0_17, n_0_16, uc_53, uc_54, uc_55, uc_56, uc_57, uc_58, 
      uc_59, uc_60, uc_61, uc_62, uc_63, uc_64, uc_65, uc_66, uc_67, uc_68, 
      uc_69}));
   datapath__0_6 i_0_5 (.p_0({n_0_719, n_0_718, n_0_717, n_0_716, n_0_715, 
      n_0_714, n_0_713, n_0_712, n_0_711, n_0_710, n_0_709, n_0_708, n_0_707, 
      n_0_706, n_0_705, multiplicand[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
      .p_1({uc_70, n_0_689, n_0_688, n_0_687, n_0_686, n_0_685, n_0_684, n_0_683, 
      n_0_682, n_0_681, n_0_680, n_0_679, n_0_678, n_0_677, n_0_676, n_0_675, 
      uc_71, uc_72, uc_73, uc_74, uc_75, uc_76, uc_77, uc_78, uc_79, uc_80, 
      uc_81, uc_82, uc_83, uc_84, uc_85, uc_86, uc_87}), .p_2({n_0_47, n_0_46, 
      n_0_45, n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, n_0_39, n_0_38, n_0_37, 
      n_0_36, n_0_35, n_0_34, n_0_33, n_0_32, uc_88, uc_89, uc_90, uc_91, uc_92, 
      uc_93, uc_94, uc_95, uc_96, uc_97, uc_98, uc_99, uc_100, uc_101, uc_102, 
      uc_103, uc_104}));
   datapath__0_7 i_0_6 (.p_0({multiplicand[15], multiplicand[14], 
      multiplicand[13], multiplicand[12], multiplicand[11], multiplicand[10], 
      multiplicand[9], multiplicand[8], multiplicand[7], multiplicand[6], 
      multiplicand[5], multiplicand[4], multiplicand[3], multiplicand[2], 
      multiplicand[1], multiplicand[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .p_1({uc_105, 
      n_0_689, n_0_688, n_0_687, n_0_686, n_0_685, n_0_684, n_0_683, n_0_682, 
      n_0_681, n_0_680, n_0_679, n_0_678, n_0_677, n_0_676, n_0_675, uc_106, 
      uc_107, uc_108, uc_109, uc_110, uc_111, uc_112, uc_113, uc_114, uc_115, 
      uc_116, uc_117, uc_118, uc_119, uc_120, uc_121, uc_122}), .p_2({n_0_63, 
      n_0_62, n_0_61, n_0_60, n_0_59, n_0_58, n_0_57, n_0_56, n_0_55, n_0_54, 
      n_0_53, n_0_52, n_0_51, n_0_50, n_0_49, n_0_48, uc_123, uc_124, uc_125, 
      uc_126, uc_127, uc_128, uc_129, uc_130, uc_131, uc_132, uc_133, uc_134, 
      uc_135, uc_136, uc_137, uc_138, uc_139}));
   datapath__0_10 i_0_8 (.p_0({n_0_719, n_0_718, n_0_717, n_0_716, n_0_715, 
      n_0_714, n_0_713, n_0_712, n_0_711, n_0_710, n_0_709, n_0_708, n_0_707, 
      n_0_706, n_0_705, multiplicand[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
      .p_1({uc_140, n_0_674, n_0_673, n_0_672, n_0_671, n_0_670, n_0_669, 
      n_0_668, n_0_667, n_0_666, n_0_665, n_0_664, n_0_663, n_0_662, n_0_661, 
      n_0_660, uc_141, uc_142, uc_143, uc_144, uc_145, uc_146, uc_147, uc_148, 
      uc_149, uc_150, uc_151, uc_152, uc_153, uc_154, uc_155, uc_156, uc_157}), 
      .p_2({n_0_79, n_0_78, n_0_77, n_0_76, n_0_75, n_0_74, n_0_73, n_0_72, 
      n_0_71, n_0_70, n_0_69, n_0_68, n_0_67, n_0_66, n_0_65, n_0_64, uc_158, 
      uc_159, uc_160, uc_161, uc_162, uc_163, uc_164, uc_165, uc_166, uc_167, 
      uc_168, uc_169, uc_170, uc_171, uc_172, uc_173, uc_174}));
   datapath__0_11 i_0_9 (.p_0({multiplicand[15], multiplicand[14], 
      multiplicand[13], multiplicand[12], multiplicand[11], multiplicand[10], 
      multiplicand[9], multiplicand[8], multiplicand[7], multiplicand[6], 
      multiplicand[5], multiplicand[4], multiplicand[3], multiplicand[2], 
      multiplicand[1], multiplicand[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .p_1({uc_175, 
      n_0_674, n_0_673, n_0_672, n_0_671, n_0_670, n_0_669, n_0_668, n_0_667, 
      n_0_666, n_0_665, n_0_664, n_0_663, n_0_662, n_0_661, n_0_660, uc_176, 
      uc_177, uc_178, uc_179, uc_180, uc_181, uc_182, uc_183, uc_184, uc_185, 
      uc_186, uc_187, uc_188, uc_189, uc_190, uc_191, uc_192}), .p_2({n_0_95, 
      n_0_94, n_0_93, n_0_92, n_0_91, n_0_90, n_0_89, n_0_88, n_0_87, n_0_86, 
      n_0_85, n_0_84, n_0_83, n_0_82, n_0_81, n_0_80, uc_193, uc_194, uc_195, 
      uc_196, uc_197, uc_198, uc_199, uc_200, uc_201, uc_202, uc_203, uc_204, 
      uc_205, uc_206, uc_207, uc_208, uc_209}));
   datapath__0_14 i_0_11 (.p_0({n_0_719, n_0_718, n_0_717, n_0_716, n_0_715, 
      n_0_714, n_0_713, n_0_712, n_0_711, n_0_710, n_0_709, n_0_708, n_0_707, 
      n_0_706, n_0_705, multiplicand[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
      .p_1({uc_210, n_0_659, n_0_658, n_0_657, n_0_656, n_0_655, n_0_654, 
      n_0_653, n_0_652, n_0_651, n_0_650, n_0_649, n_0_648, n_0_647, n_0_646, 
      n_0_645, uc_211, uc_212, uc_213, uc_214, uc_215, uc_216, uc_217, uc_218, 
      uc_219, uc_220, uc_221, uc_222, uc_223, uc_224, uc_225, uc_226, uc_227}), 
      .p_2({n_0_111, n_0_110, n_0_109, n_0_108, n_0_107, n_0_106, n_0_105, 
      n_0_104, n_0_103, n_0_102, n_0_101, n_0_100, n_0_99, n_0_98, n_0_97, 
      n_0_96, uc_228, uc_229, uc_230, uc_231, uc_232, uc_233, uc_234, uc_235, 
      uc_236, uc_237, uc_238, uc_239, uc_240, uc_241, uc_242, uc_243, uc_244}));
   datapath__0_15 i_0_12 (.p_0({multiplicand[15], multiplicand[14], 
      multiplicand[13], multiplicand[12], multiplicand[11], multiplicand[10], 
      multiplicand[9], multiplicand[8], multiplicand[7], multiplicand[6], 
      multiplicand[5], multiplicand[4], multiplicand[3], multiplicand[2], 
      multiplicand[1], multiplicand[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .p_1({uc_245, 
      n_0_659, n_0_658, n_0_657, n_0_656, n_0_655, n_0_654, n_0_653, n_0_652, 
      n_0_651, n_0_650, n_0_649, n_0_648, n_0_647, n_0_646, n_0_645, uc_246, 
      uc_247, uc_248, uc_249, uc_250, uc_251, uc_252, uc_253, uc_254, uc_255, 
      uc_256, uc_257, uc_258, uc_259, uc_260, uc_261, uc_262}), .p_2({n_0_127, 
      n_0_126, n_0_125, n_0_124, n_0_123, n_0_122, n_0_121, n_0_120, n_0_119, 
      n_0_118, n_0_117, n_0_116, n_0_115, n_0_114, n_0_113, n_0_112, uc_263, 
      uc_264, uc_265, uc_266, uc_267, uc_268, uc_269, uc_270, uc_271, uc_272, 
      uc_273, uc_274, uc_275, uc_276, uc_277, uc_278, uc_279}));
   datapath__0_18 i_0_14 (.p_0({n_0_719, n_0_718, n_0_717, n_0_716, n_0_715, 
      n_0_714, n_0_713, n_0_712, n_0_711, n_0_710, n_0_709, n_0_708, n_0_707, 
      n_0_706, n_0_705, multiplicand[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
      .p_1({uc_280, n_0_644, n_0_643, n_0_642, n_0_641, n_0_640, n_0_639, 
      n_0_638, n_0_637, n_0_636, n_0_635, n_0_634, n_0_633, n_0_632, n_0_631, 
      n_0_630, uc_281, uc_282, uc_283, uc_284, uc_285, uc_286, uc_287, uc_288, 
      uc_289, uc_290, uc_291, uc_292, uc_293, uc_294, uc_295, uc_296, uc_297}), 
      .p_2({n_0_143, n_0_142, n_0_141, n_0_140, n_0_139, n_0_138, n_0_137, 
      n_0_136, n_0_135, n_0_134, n_0_133, n_0_132, n_0_131, n_0_130, n_0_129, 
      n_0_128, uc_298, uc_299, uc_300, uc_301, uc_302, uc_303, uc_304, uc_305, 
      uc_306, uc_307, uc_308, uc_309, uc_310, uc_311, uc_312, uc_313, uc_314}));
   datapath__0_19 i_0_15 (.p_0({multiplicand[15], multiplicand[14], 
      multiplicand[13], multiplicand[12], multiplicand[11], multiplicand[10], 
      multiplicand[9], multiplicand[8], multiplicand[7], multiplicand[6], 
      multiplicand[5], multiplicand[4], multiplicand[3], multiplicand[2], 
      multiplicand[1], multiplicand[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .p_1({uc_315, 
      n_0_644, n_0_643, n_0_642, n_0_641, n_0_640, n_0_639, n_0_638, n_0_637, 
      n_0_636, n_0_635, n_0_634, n_0_633, n_0_632, n_0_631, n_0_630, uc_316, 
      uc_317, uc_318, uc_319, uc_320, uc_321, uc_322, uc_323, uc_324, uc_325, 
      uc_326, uc_327, uc_328, uc_329, uc_330, uc_331, uc_332}), .p_2({n_0_159, 
      n_0_158, n_0_157, n_0_156, n_0_155, n_0_154, n_0_153, n_0_152, n_0_151, 
      n_0_150, n_0_149, n_0_148, n_0_147, n_0_146, n_0_145, n_0_144, uc_333, 
      uc_334, uc_335, uc_336, uc_337, uc_338, uc_339, uc_340, uc_341, uc_342, 
      uc_343, uc_344, uc_345, uc_346, uc_347, uc_348, uc_349}));
   datapath__0_22 i_0_17 (.p_0({n_0_719, n_0_718, n_0_717, n_0_716, n_0_715, 
      n_0_714, n_0_713, n_0_712, n_0_711, n_0_710, n_0_709, n_0_708, n_0_707, 
      n_0_706, n_0_705, multiplicand[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
      .p_1({uc_350, n_0_629, n_0_628, n_0_627, n_0_626, n_0_625, n_0_624, 
      n_0_623, n_0_622, n_0_621, n_0_620, n_0_619, n_0_618, n_0_617, n_0_616, 
      n_0_615, uc_351, uc_352, uc_353, uc_354, uc_355, uc_356, uc_357, uc_358, 
      uc_359, uc_360, uc_361, uc_362, uc_363, uc_364, uc_365, uc_366, uc_367}), 
      .p_2({n_0_175, n_0_174, n_0_173, n_0_172, n_0_171, n_0_170, n_0_169, 
      n_0_168, n_0_167, n_0_166, n_0_165, n_0_164, n_0_163, n_0_162, n_0_161, 
      n_0_160, uc_368, uc_369, uc_370, uc_371, uc_372, uc_373, uc_374, uc_375, 
      uc_376, uc_377, uc_378, uc_379, uc_380, uc_381, uc_382, uc_383, uc_384}));
   datapath__0_23 i_0_18 (.p_0({multiplicand[15], multiplicand[14], 
      multiplicand[13], multiplicand[12], multiplicand[11], multiplicand[10], 
      multiplicand[9], multiplicand[8], multiplicand[7], multiplicand[6], 
      multiplicand[5], multiplicand[4], multiplicand[3], multiplicand[2], 
      multiplicand[1], multiplicand[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .p_1({uc_385, 
      n_0_629, n_0_628, n_0_627, n_0_626, n_0_625, n_0_624, n_0_623, n_0_622, 
      n_0_621, n_0_620, n_0_619, n_0_618, n_0_617, n_0_616, n_0_615, uc_386, 
      uc_387, uc_388, uc_389, uc_390, uc_391, uc_392, uc_393, uc_394, uc_395, 
      uc_396, uc_397, uc_398, uc_399, uc_400, uc_401, uc_402}), .p_2({n_0_191, 
      n_0_190, n_0_189, n_0_188, n_0_187, n_0_186, n_0_185, n_0_184, n_0_183, 
      n_0_182, n_0_181, n_0_180, n_0_179, n_0_178, n_0_177, n_0_176, uc_403, 
      uc_404, uc_405, uc_406, uc_407, uc_408, uc_409, uc_410, uc_411, uc_412, 
      uc_413, uc_414, uc_415, uc_416, uc_417, uc_418, uc_419}));
   datapath__0_26 i_0_20 (.p_0({n_0_719, n_0_718, n_0_717, n_0_716, n_0_715, 
      n_0_714, n_0_713, n_0_712, n_0_711, n_0_710, n_0_709, n_0_708, n_0_707, 
      n_0_706, n_0_705, multiplicand[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
      .p_1({uc_420, n_0_614, n_0_613, n_0_612, n_0_611, n_0_610, n_0_609, 
      n_0_608, n_0_607, n_0_606, n_0_605, n_0_604, n_0_603, n_0_602, n_0_601, 
      n_0_600, uc_421, uc_422, uc_423, uc_424, uc_425, uc_426, uc_427, uc_428, 
      uc_429, uc_430, uc_431, uc_432, uc_433, uc_434, uc_435, uc_436, uc_437}), 
      .p_2({n_0_207, n_0_206, n_0_205, n_0_204, n_0_203, n_0_202, n_0_201, 
      n_0_200, n_0_199, n_0_198, n_0_197, n_0_196, n_0_195, n_0_194, n_0_193, 
      n_0_192, uc_438, uc_439, uc_440, uc_441, uc_442, uc_443, uc_444, uc_445, 
      uc_446, uc_447, uc_448, uc_449, uc_450, uc_451, uc_452, uc_453, uc_454}));
   datapath__0_27 i_0_21 (.p_0({multiplicand[15], multiplicand[14], 
      multiplicand[13], multiplicand[12], multiplicand[11], multiplicand[10], 
      multiplicand[9], multiplicand[8], multiplicand[7], multiplicand[6], 
      multiplicand[5], multiplicand[4], multiplicand[3], multiplicand[2], 
      multiplicand[1], multiplicand[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .p_1({uc_455, 
      n_0_614, n_0_613, n_0_612, n_0_611, n_0_610, n_0_609, n_0_608, n_0_607, 
      n_0_606, n_0_605, n_0_604, n_0_603, n_0_602, n_0_601, n_0_600, uc_456, 
      uc_457, uc_458, uc_459, uc_460, uc_461, uc_462, uc_463, uc_464, uc_465, 
      uc_466, uc_467, uc_468, uc_469, uc_470, uc_471, uc_472}), .p_2({n_0_223, 
      n_0_222, n_0_221, n_0_220, n_0_219, n_0_218, n_0_217, n_0_216, n_0_215, 
      n_0_214, n_0_213, n_0_212, n_0_211, n_0_210, n_0_209, n_0_208, uc_473, 
      uc_474, uc_475, uc_476, uc_477, uc_478, uc_479, uc_480, uc_481, uc_482, 
      uc_483, uc_484, uc_485, uc_486, uc_487, uc_488, uc_489}));
   datapath__0_30 i_0_23 (.p_0({n_0_719, n_0_718, n_0_717, n_0_716, n_0_715, 
      n_0_714, n_0_713, n_0_712, n_0_711, n_0_710, n_0_709, n_0_708, n_0_707, 
      n_0_706, n_0_705, multiplicand[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
      .p_1({uc_490, n_0_599, n_0_598, n_0_597, n_0_596, n_0_595, n_0_594, 
      n_0_593, n_0_592, n_0_591, n_0_590, n_0_589, n_0_588, n_0_587, n_0_586, 
      n_0_585, uc_491, uc_492, uc_493, uc_494, uc_495, uc_496, uc_497, uc_498, 
      uc_499, uc_500, uc_501, uc_502, uc_503, uc_504, uc_505, uc_506, uc_507}), 
      .p_2({n_0_239, n_0_238, n_0_237, n_0_236, n_0_235, n_0_234, n_0_233, 
      n_0_232, n_0_231, n_0_230, n_0_229, n_0_228, n_0_227, n_0_226, n_0_225, 
      n_0_224, uc_508, uc_509, uc_510, uc_511, uc_512, uc_513, uc_514, uc_515, 
      uc_516, uc_517, uc_518, uc_519, uc_520, uc_521, uc_522, uc_523, uc_524}));
   datapath__0_31 i_0_24 (.p_0({multiplicand[15], multiplicand[14], 
      multiplicand[13], multiplicand[12], multiplicand[11], multiplicand[10], 
      multiplicand[9], multiplicand[8], multiplicand[7], multiplicand[6], 
      multiplicand[5], multiplicand[4], multiplicand[3], multiplicand[2], 
      multiplicand[1], multiplicand[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .p_1({uc_525, 
      n_0_599, n_0_598, n_0_597, n_0_596, n_0_595, n_0_594, n_0_593, n_0_592, 
      n_0_591, n_0_590, n_0_589, n_0_588, n_0_587, n_0_586, n_0_585, uc_526, 
      uc_527, uc_528, uc_529, uc_530, uc_531, uc_532, uc_533, uc_534, uc_535, 
      uc_536, uc_537, uc_538, uc_539, uc_540, uc_541, uc_542}), .p_2({n_0_255, 
      n_0_254, n_0_253, n_0_252, n_0_251, n_0_250, n_0_249, n_0_248, n_0_247, 
      n_0_246, n_0_245, n_0_244, n_0_243, n_0_242, n_0_241, n_0_240, uc_543, 
      uc_544, uc_545, uc_546, uc_547, uc_548, uc_549, uc_550, uc_551, uc_552, 
      uc_553, uc_554, uc_555, uc_556, uc_557, uc_558, uc_559}));
   datapath__0_34 i_0_26 (.p_0({n_0_719, n_0_718, n_0_717, n_0_716, n_0_715, 
      n_0_714, n_0_713, n_0_712, n_0_711, n_0_710, n_0_709, n_0_708, n_0_707, 
      n_0_706, n_0_705, multiplicand[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
      .p_1({uc_560, n_0_584, n_0_583, n_0_582, n_0_581, n_0_580, n_0_579, 
      n_0_578, n_0_577, n_0_576, n_0_575, n_0_574, n_0_573, n_0_572, n_0_571, 
      n_0_570, uc_561, uc_562, uc_563, uc_564, uc_565, uc_566, uc_567, uc_568, 
      uc_569, uc_570, uc_571, uc_572, uc_573, uc_574, uc_575, uc_576, uc_577}), 
      .p_2({n_0_271, n_0_270, n_0_269, n_0_268, n_0_267, n_0_266, n_0_265, 
      n_0_264, n_0_263, n_0_262, n_0_261, n_0_260, n_0_259, n_0_258, n_0_257, 
      n_0_256, uc_578, uc_579, uc_580, uc_581, uc_582, uc_583, uc_584, uc_585, 
      uc_586, uc_587, uc_588, uc_589, uc_590, uc_591, uc_592, uc_593, uc_594}));
   datapath__0_35 i_0_27 (.p_0({multiplicand[15], multiplicand[14], 
      multiplicand[13], multiplicand[12], multiplicand[11], multiplicand[10], 
      multiplicand[9], multiplicand[8], multiplicand[7], multiplicand[6], 
      multiplicand[5], multiplicand[4], multiplicand[3], multiplicand[2], 
      multiplicand[1], multiplicand[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .p_1({uc_595, 
      n_0_584, n_0_583, n_0_582, n_0_581, n_0_580, n_0_579, n_0_578, n_0_577, 
      n_0_576, n_0_575, n_0_574, n_0_573, n_0_572, n_0_571, n_0_570, uc_596, 
      uc_597, uc_598, uc_599, uc_600, uc_601, uc_602, uc_603, uc_604, uc_605, 
      uc_606, uc_607, uc_608, uc_609, uc_610, uc_611, uc_612}), .p_2({n_0_287, 
      n_0_286, n_0_285, n_0_284, n_0_283, n_0_282, n_0_281, n_0_280, n_0_279, 
      n_0_278, n_0_277, n_0_276, n_0_275, n_0_274, n_0_273, n_0_272, uc_613, 
      uc_614, uc_615, uc_616, uc_617, uc_618, uc_619, uc_620, uc_621, uc_622, 
      uc_623, uc_624, uc_625, uc_626, uc_627, uc_628, uc_629}));
   datapath__0_38 i_0_29 (.p_0({n_0_719, n_0_718, n_0_717, n_0_716, n_0_715, 
      n_0_714, n_0_713, n_0_712, n_0_711, n_0_710, n_0_709, n_0_708, n_0_707, 
      n_0_706, n_0_705, multiplicand[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
      .p_1({uc_630, n_0_569, n_0_568, n_0_567, n_0_566, n_0_565, n_0_564, 
      n_0_563, n_0_562, n_0_561, n_0_560, n_0_559, n_0_558, n_0_557, n_0_556, 
      n_0_555, uc_631, uc_632, uc_633, uc_634, uc_635, uc_636, uc_637, uc_638, 
      uc_639, uc_640, uc_641, uc_642, uc_643, uc_644, uc_645, uc_646, uc_647}), 
      .p_2({n_0_303, n_0_302, n_0_301, n_0_300, n_0_299, n_0_298, n_0_297, 
      n_0_296, n_0_295, n_0_294, n_0_293, n_0_292, n_0_291, n_0_290, n_0_289, 
      n_0_288, uc_648, uc_649, uc_650, uc_651, uc_652, uc_653, uc_654, uc_655, 
      uc_656, uc_657, uc_658, uc_659, uc_660, uc_661, uc_662, uc_663, uc_664}));
   datapath__0_39 i_0_30 (.p_0({multiplicand[15], multiplicand[14], 
      multiplicand[13], multiplicand[12], multiplicand[11], multiplicand[10], 
      multiplicand[9], multiplicand[8], multiplicand[7], multiplicand[6], 
      multiplicand[5], multiplicand[4], multiplicand[3], multiplicand[2], 
      multiplicand[1], multiplicand[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .p_1({uc_665, 
      n_0_569, n_0_568, n_0_567, n_0_566, n_0_565, n_0_564, n_0_563, n_0_562, 
      n_0_561, n_0_560, n_0_559, n_0_558, n_0_557, n_0_556, n_0_555, uc_666, 
      uc_667, uc_668, uc_669, uc_670, uc_671, uc_672, uc_673, uc_674, uc_675, 
      uc_676, uc_677, uc_678, uc_679, uc_680, uc_681, uc_682}), .p_2({n_0_319, 
      n_0_318, n_0_317, n_0_316, n_0_315, n_0_314, n_0_313, n_0_312, n_0_311, 
      n_0_310, n_0_309, n_0_308, n_0_307, n_0_306, n_0_305, n_0_304, uc_683, 
      uc_684, uc_685, uc_686, uc_687, uc_688, uc_689, uc_690, uc_691, uc_692, 
      uc_693, uc_694, uc_695, uc_696, uc_697, uc_698, uc_699}));
   datapath__0_42 i_0_32 (.p_0({n_0_719, n_0_718, n_0_717, n_0_716, n_0_715, 
      n_0_714, n_0_713, n_0_712, n_0_711, n_0_710, n_0_709, n_0_708, n_0_707, 
      n_0_706, n_0_705, multiplicand[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
      .p_1({uc_700, n_0_554, n_0_553, n_0_552, n_0_551, n_0_550, n_0_549, 
      n_0_548, n_0_547, n_0_546, n_0_545, n_0_544, n_0_543, n_0_542, n_0_541, 
      n_0_540, uc_701, uc_702, uc_703, uc_704, uc_705, uc_706, uc_707, uc_708, 
      uc_709, uc_710, uc_711, uc_712, uc_713, uc_714, uc_715, uc_716, uc_717}), 
      .p_2({n_0_335, n_0_334, n_0_333, n_0_332, n_0_331, n_0_330, n_0_329, 
      n_0_328, n_0_327, n_0_326, n_0_325, n_0_324, n_0_323, n_0_322, n_0_321, 
      n_0_320, uc_718, uc_719, uc_720, uc_721, uc_722, uc_723, uc_724, uc_725, 
      uc_726, uc_727, uc_728, uc_729, uc_730, uc_731, uc_732, uc_733, uc_734}));
   datapath__0_43 i_0_33 (.p_0({multiplicand[15], multiplicand[14], 
      multiplicand[13], multiplicand[12], multiplicand[11], multiplicand[10], 
      multiplicand[9], multiplicand[8], multiplicand[7], multiplicand[6], 
      multiplicand[5], multiplicand[4], multiplicand[3], multiplicand[2], 
      multiplicand[1], multiplicand[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .p_1({uc_735, 
      n_0_554, n_0_553, n_0_552, n_0_551, n_0_550, n_0_549, n_0_548, n_0_547, 
      n_0_546, n_0_545, n_0_544, n_0_543, n_0_542, n_0_541, n_0_540, uc_736, 
      uc_737, uc_738, uc_739, uc_740, uc_741, uc_742, uc_743, uc_744, uc_745, 
      uc_746, uc_747, uc_748, uc_749, uc_750, uc_751, uc_752}), .p_2({n_0_351, 
      n_0_350, n_0_349, n_0_348, n_0_347, n_0_346, n_0_345, n_0_344, n_0_343, 
      n_0_342, n_0_341, n_0_340, n_0_339, n_0_338, n_0_337, n_0_336, uc_753, 
      uc_754, uc_755, uc_756, uc_757, uc_758, uc_759, uc_760, uc_761, uc_762, 
      uc_763, uc_764, uc_765, uc_766, uc_767, uc_768, uc_769}));
   datapath__0_46 i_0_35 (.p_0({n_0_719, n_0_718, n_0_717, n_0_716, n_0_715, 
      n_0_714, n_0_713, n_0_712, n_0_711, n_0_710, n_0_709, n_0_708, n_0_707, 
      n_0_706, n_0_705, multiplicand[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
      .p_1({uc_770, n_0_539, n_0_538, n_0_537, n_0_536, n_0_535, n_0_534, 
      n_0_533, n_0_532, n_0_531, n_0_530, n_0_529, n_0_528, n_0_527, n_0_526, 
      n_0_525, uc_771, uc_772, uc_773, uc_774, uc_775, uc_776, uc_777, uc_778, 
      uc_779, uc_780, uc_781, uc_782, uc_783, uc_784, uc_785, uc_786, uc_787}), 
      .p_2({n_0_367, n_0_366, n_0_365, n_0_364, n_0_363, n_0_362, n_0_361, 
      n_0_360, n_0_359, n_0_358, n_0_357, n_0_356, n_0_355, n_0_354, n_0_353, 
      n_0_352, uc_788, uc_789, uc_790, uc_791, uc_792, uc_793, uc_794, uc_795, 
      uc_796, uc_797, uc_798, uc_799, uc_800, uc_801, uc_802, uc_803, uc_804}));
   datapath__0_47 i_0_36 (.p_0({multiplicand[15], multiplicand[14], 
      multiplicand[13], multiplicand[12], multiplicand[11], multiplicand[10], 
      multiplicand[9], multiplicand[8], multiplicand[7], multiplicand[6], 
      multiplicand[5], multiplicand[4], multiplicand[3], multiplicand[2], 
      multiplicand[1], multiplicand[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .p_1({uc_805, 
      n_0_539, n_0_538, n_0_537, n_0_536, n_0_535, n_0_534, n_0_533, n_0_532, 
      n_0_531, n_0_530, n_0_529, n_0_528, n_0_527, n_0_526, n_0_525, uc_806, 
      uc_807, uc_808, uc_809, uc_810, uc_811, uc_812, uc_813, uc_814, uc_815, 
      uc_816, uc_817, uc_818, uc_819, uc_820, uc_821, uc_822}), .p_2({n_0_383, 
      n_0_382, n_0_381, n_0_380, n_0_379, n_0_378, n_0_377, n_0_376, n_0_375, 
      n_0_374, n_0_373, n_0_372, n_0_371, n_0_370, n_0_369, n_0_368, uc_823, 
      uc_824, uc_825, uc_826, uc_827, uc_828, uc_829, uc_830, uc_831, uc_832, 
      uc_833, uc_834, uc_835, uc_836, uc_837, uc_838, uc_839}));
   datapath__0_50 i_0_38 (.p_0({n_0_719, n_0_718, n_0_717, n_0_716, n_0_715, 
      n_0_714, n_0_713, n_0_712, n_0_711, n_0_710, n_0_709, n_0_708, n_0_707, 
      n_0_706, n_0_705, multiplicand[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
      .p_1({uc_840, n_0_524, n_0_523, n_0_522, n_0_521, n_0_520, n_0_519, 
      n_0_518, n_0_517, n_0_516, n_0_515, n_0_514, n_0_513, n_0_512, n_0_511, 
      n_0_510, uc_841, uc_842, uc_843, uc_844, uc_845, uc_846, uc_847, uc_848, 
      uc_849, uc_850, uc_851, uc_852, uc_853, uc_854, uc_855, uc_856, uc_857}), 
      .p_2({n_0_399, n_0_398, n_0_397, n_0_396, n_0_395, n_0_394, n_0_393, 
      n_0_392, n_0_391, n_0_390, n_0_389, n_0_388, n_0_387, n_0_386, n_0_385, 
      n_0_384, uc_858, uc_859, uc_860, uc_861, uc_862, uc_863, uc_864, uc_865, 
      uc_866, uc_867, uc_868, uc_869, uc_870, uc_871, uc_872, uc_873, uc_874}));
   datapath__0_51 i_0_39 (.p_0({multiplicand[15], multiplicand[14], 
      multiplicand[13], multiplicand[12], multiplicand[11], multiplicand[10], 
      multiplicand[9], multiplicand[8], multiplicand[7], multiplicand[6], 
      multiplicand[5], multiplicand[4], multiplicand[3], multiplicand[2], 
      multiplicand[1], multiplicand[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .p_1({uc_875, 
      n_0_524, n_0_523, n_0_522, n_0_521, n_0_520, n_0_519, n_0_518, n_0_517, 
      n_0_516, n_0_515, n_0_514, n_0_513, n_0_512, n_0_511, n_0_510, uc_876, 
      uc_877, uc_878, uc_879, uc_880, uc_881, uc_882, uc_883, uc_884, uc_885, 
      uc_886, uc_887, uc_888, uc_889, uc_890, uc_891, uc_892}), .p_2({n_0_415, 
      n_0_414, n_0_413, n_0_412, n_0_411, n_0_410, n_0_409, n_0_408, n_0_407, 
      n_0_406, n_0_405, n_0_404, n_0_403, n_0_402, n_0_401, n_0_400, uc_893, 
      uc_894, uc_895, uc_896, uc_897, uc_898, uc_899, uc_900, uc_901, uc_902, 
      uc_903, uc_904, uc_905, uc_906, uc_907, uc_908, uc_909}));
   datapath__0_54 i_0_41 (.p_0({n_0_719, n_0_718, n_0_717, n_0_716, n_0_715, 
      n_0_714, n_0_713, n_0_712, n_0_711, n_0_710, n_0_709, n_0_708, n_0_707, 
      n_0_706, n_0_705, multiplicand[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
      .p_1({uc_910, n_0_509, n_0_508, n_0_507, n_0_506, n_0_505, n_0_504, 
      n_0_503, n_0_502, n_0_501, n_0_500, n_0_499, n_0_498, n_0_497, n_0_496, 
      n_0_495, uc_911, uc_912, uc_913, uc_914, uc_915, uc_916, uc_917, uc_918, 
      uc_919, uc_920, uc_921, uc_922, uc_923, uc_924, uc_925, uc_926, uc_927}), 
      .p_2({n_0_431, n_0_430, n_0_429, n_0_428, n_0_427, n_0_426, n_0_425, 
      n_0_424, n_0_423, n_0_422, n_0_421, n_0_420, n_0_419, n_0_418, n_0_417, 
      n_0_416, uc_928, uc_929, uc_930, uc_931, uc_932, uc_933, uc_934, uc_935, 
      uc_936, uc_937, uc_938, uc_939, uc_940, uc_941, uc_942, uc_943, uc_944}));
   datapath__0_55 i_0_42 (.p_0({multiplicand[15], multiplicand[14], 
      multiplicand[13], multiplicand[12], multiplicand[11], multiplicand[10], 
      multiplicand[9], multiplicand[8], multiplicand[7], multiplicand[6], 
      multiplicand[5], multiplicand[4], multiplicand[3], multiplicand[2], 
      multiplicand[1], multiplicand[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .p_1({uc_945, 
      n_0_509, n_0_508, n_0_507, n_0_506, n_0_505, n_0_504, n_0_503, n_0_502, 
      n_0_501, n_0_500, n_0_499, n_0_498, n_0_497, n_0_496, n_0_495, uc_946, 
      uc_947, uc_948, uc_949, uc_950, uc_951, uc_952, uc_953, uc_954, uc_955, 
      uc_956, uc_957, uc_958, uc_959, uc_960, uc_961, uc_962}), .p_2({n_0_447, 
      n_0_446, n_0_445, n_0_444, n_0_443, n_0_442, n_0_441, n_0_440, n_0_439, 
      n_0_438, n_0_437, n_0_436, n_0_435, n_0_434, n_0_433, n_0_432, uc_963, 
      uc_964, uc_965, uc_966, uc_967, uc_968, uc_969, uc_970, uc_971, uc_972, 
      uc_973, uc_974, uc_975, uc_976, uc_977, uc_978, uc_979}));
   datapath__0_58 i_0_44 (.p_0({n_0_719, n_0_718, n_0_717, n_0_716, n_0_715, 
      n_0_714, n_0_713, n_0_712, n_0_711, n_0_710, n_0_709, n_0_708, n_0_707, 
      n_0_706, n_0_705, multiplicand[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
      .p_1({uc_980, n_0_494, n_0_493, n_0_492, n_0_491, n_0_490, n_0_489, 
      n_0_488, n_0_487, n_0_486, n_0_485, n_0_484, n_0_483, n_0_482, n_0_481, 
      n_0_480, uc_981, uc_982, uc_983, uc_984, uc_985, uc_986, uc_987, uc_988, 
      uc_989, uc_990, uc_991, uc_992, uc_993, uc_994, uc_995, uc_996, uc_997}), 
      .p_2({n_0_463, n_0_462, n_0_461, n_0_460, n_0_459, n_0_458, n_0_457, 
      n_0_456, n_0_455, n_0_454, n_0_453, n_0_452, n_0_451, n_0_450, n_0_449, 
      n_0_448, uc_998, uc_999, uc_1000, uc_1001, uc_1002, uc_1003, uc_1004, 
      uc_1005, uc_1006, uc_1007, uc_1008, uc_1009, uc_1010, uc_1011, uc_1012, 
      uc_1013, uc_1014}));
   datapath__0_59 i_0_45 (.p_0({multiplicand[15], multiplicand[14], 
      multiplicand[13], multiplicand[12], multiplicand[11], multiplicand[10], 
      multiplicand[9], multiplicand[8], multiplicand[7], multiplicand[6], 
      multiplicand[5], multiplicand[4], multiplicand[3], multiplicand[2], 
      multiplicand[1], multiplicand[0], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .p_1({
      uc_1015, n_0_494, n_0_493, n_0_492, n_0_491, n_0_490, n_0_489, n_0_488, 
      n_0_487, n_0_486, n_0_485, n_0_484, n_0_483, n_0_482, n_0_481, n_0_480, 
      uc_1016, uc_1017, uc_1018, uc_1019, uc_1020, uc_1021, uc_1022, uc_1023, 
      uc_1024, uc_1025, uc_1026, uc_1027, uc_1028, uc_1029, uc_1030, uc_1031, 
      uc_1032}), .p_2({n_0_479, n_0_478, n_0_477, n_0_476, n_0_475, n_0_474, 
      n_0_473, n_0_472, n_0_471, n_0_470, n_0_469, n_0_468, n_0_467, n_0_466, 
      n_0_465, n_0_464, uc_1033, uc_1034, uc_1035, uc_1036, uc_1037, uc_1038, 
      uc_1039, uc_1040, uc_1041, uc_1042, uc_1043, uc_1044, uc_1045, uc_1046, 
      uc_1047, uc_1048, uc_1049}));
   INV_X1 i_0_0_0 (.A(n_0_0_0), .ZN(product[15]));
   AOI222_X1 i_0_0_1 (.A1(n_0_448), .A2(n_0_0_19), .B1(n_0_464), .B2(n_0_0_18), 
      .C1(n_0_480), .C2(n_0_0_17), .ZN(n_0_0_0));
   INV_X1 i_0_0_2 (.A(n_0_0_1), .ZN(product[16]));
   AOI222_X1 i_0_0_3 (.A1(n_0_449), .A2(n_0_0_19), .B1(n_0_465), .B2(n_0_0_18), 
      .C1(n_0_481), .C2(n_0_0_17), .ZN(n_0_0_1));
   INV_X1 i_0_0_4 (.A(n_0_0_2), .ZN(product[17]));
   AOI222_X1 i_0_0_5 (.A1(n_0_450), .A2(n_0_0_19), .B1(n_0_466), .B2(n_0_0_18), 
      .C1(n_0_482), .C2(n_0_0_17), .ZN(n_0_0_2));
   INV_X1 i_0_0_6 (.A(n_0_0_3), .ZN(product[18]));
   AOI222_X1 i_0_0_7 (.A1(n_0_451), .A2(n_0_0_19), .B1(n_0_467), .B2(n_0_0_18), 
      .C1(n_0_483), .C2(n_0_0_17), .ZN(n_0_0_3));
   INV_X1 i_0_0_8 (.A(n_0_0_4), .ZN(product[19]));
   AOI222_X1 i_0_0_9 (.A1(n_0_452), .A2(n_0_0_19), .B1(n_0_468), .B2(n_0_0_18), 
      .C1(n_0_484), .C2(n_0_0_17), .ZN(n_0_0_4));
   INV_X1 i_0_0_10 (.A(n_0_0_5), .ZN(product[20]));
   AOI222_X1 i_0_0_11 (.A1(n_0_453), .A2(n_0_0_19), .B1(n_0_469), .B2(n_0_0_18), 
      .C1(n_0_485), .C2(n_0_0_17), .ZN(n_0_0_5));
   INV_X1 i_0_0_12 (.A(n_0_0_6), .ZN(product[21]));
   AOI222_X1 i_0_0_13 (.A1(n_0_454), .A2(n_0_0_19), .B1(n_0_470), .B2(n_0_0_18), 
      .C1(n_0_486), .C2(n_0_0_17), .ZN(n_0_0_6));
   INV_X1 i_0_0_14 (.A(n_0_0_7), .ZN(product[22]));
   AOI222_X1 i_0_0_15 (.A1(n_0_455), .A2(n_0_0_19), .B1(n_0_471), .B2(n_0_0_18), 
      .C1(n_0_487), .C2(n_0_0_17), .ZN(n_0_0_7));
   INV_X1 i_0_0_16 (.A(n_0_0_8), .ZN(product[23]));
   AOI222_X1 i_0_0_17 (.A1(n_0_456), .A2(n_0_0_19), .B1(n_0_472), .B2(n_0_0_18), 
      .C1(n_0_488), .C2(n_0_0_17), .ZN(n_0_0_8));
   INV_X1 i_0_0_18 (.A(n_0_0_9), .ZN(product[24]));
   AOI222_X1 i_0_0_19 (.A1(n_0_457), .A2(n_0_0_19), .B1(n_0_473), .B2(n_0_0_18), 
      .C1(n_0_489), .C2(n_0_0_17), .ZN(n_0_0_9));
   INV_X1 i_0_0_20 (.A(n_0_0_10), .ZN(product[25]));
   AOI222_X1 i_0_0_21 (.A1(n_0_458), .A2(n_0_0_19), .B1(n_0_474), .B2(n_0_0_18), 
      .C1(n_0_490), .C2(n_0_0_17), .ZN(n_0_0_10));
   INV_X1 i_0_0_22 (.A(n_0_0_11), .ZN(product[26]));
   AOI222_X1 i_0_0_23 (.A1(n_0_459), .A2(n_0_0_19), .B1(n_0_475), .B2(n_0_0_18), 
      .C1(n_0_491), .C2(n_0_0_17), .ZN(n_0_0_11));
   INV_X1 i_0_0_24 (.A(n_0_0_12), .ZN(product[27]));
   AOI222_X1 i_0_0_25 (.A1(n_0_460), .A2(n_0_0_19), .B1(n_0_476), .B2(n_0_0_18), 
      .C1(n_0_492), .C2(n_0_0_17), .ZN(n_0_0_12));
   INV_X1 i_0_0_26 (.A(n_0_0_13), .ZN(product[28]));
   AOI222_X1 i_0_0_27 (.A1(n_0_461), .A2(n_0_0_19), .B1(n_0_477), .B2(n_0_0_18), 
      .C1(n_0_493), .C2(n_0_0_17), .ZN(n_0_0_13));
   INV_X1 i_0_0_28 (.A(n_0_0_14), .ZN(product[29]));
   AOI221_X1 i_0_0_29 (.A(n_0_0_16), .B1(n_0_462), .B2(n_0_0_19), .C1(n_0_478), 
      .C2(n_0_0_18), .ZN(n_0_0_14));
   INV_X1 i_0_0_30 (.A(n_0_0_15), .ZN(product[30]));
   AOI221_X1 i_0_0_31 (.A(n_0_0_16), .B1(n_0_463), .B2(n_0_0_19), .C1(n_0_479), 
      .C2(n_0_0_18), .ZN(n_0_0_15));
   AND2_X1 i_0_0_32 (.A1(n_0_494), .A2(n_0_0_17), .ZN(n_0_0_16));
   NOR2_X1 i_0_0_33 (.A1(n_0_0_19), .A2(n_0_0_18), .ZN(n_0_0_17));
   NOR2_X1 i_0_0_34 (.A1(multiplier[15]), .A2(n_0_0_341), .ZN(n_0_0_18));
   AND2_X1 i_0_0_35 (.A1(multiplier[15]), .A2(n_0_0_341), .ZN(n_0_0_19));
   INV_X1 i_0_0_36 (.A(n_0_0_20), .ZN(product[14]));
   AOI222_X1 i_0_0_37 (.A1(n_0_416), .A2(n_0_0_39), .B1(n_0_432), .B2(n_0_0_38), 
      .C1(n_0_495), .C2(n_0_0_37), .ZN(n_0_0_20));
   INV_X1 i_0_0_38 (.A(n_0_0_21), .ZN(n_0_480));
   AOI222_X1 i_0_0_39 (.A1(n_0_417), .A2(n_0_0_39), .B1(n_0_433), .B2(n_0_0_38), 
      .C1(n_0_496), .C2(n_0_0_37), .ZN(n_0_0_21));
   INV_X1 i_0_0_40 (.A(n_0_0_22), .ZN(n_0_481));
   AOI222_X1 i_0_0_41 (.A1(n_0_418), .A2(n_0_0_39), .B1(n_0_434), .B2(n_0_0_38), 
      .C1(n_0_497), .C2(n_0_0_37), .ZN(n_0_0_22));
   INV_X1 i_0_0_42 (.A(n_0_0_23), .ZN(n_0_482));
   AOI222_X1 i_0_0_43 (.A1(n_0_419), .A2(n_0_0_39), .B1(n_0_435), .B2(n_0_0_38), 
      .C1(n_0_498), .C2(n_0_0_37), .ZN(n_0_0_23));
   INV_X1 i_0_0_44 (.A(n_0_0_24), .ZN(n_0_483));
   AOI222_X1 i_0_0_45 (.A1(n_0_420), .A2(n_0_0_39), .B1(n_0_436), .B2(n_0_0_38), 
      .C1(n_0_499), .C2(n_0_0_37), .ZN(n_0_0_24));
   INV_X1 i_0_0_46 (.A(n_0_0_25), .ZN(n_0_484));
   AOI222_X1 i_0_0_47 (.A1(n_0_421), .A2(n_0_0_39), .B1(n_0_437), .B2(n_0_0_38), 
      .C1(n_0_500), .C2(n_0_0_37), .ZN(n_0_0_25));
   INV_X1 i_0_0_48 (.A(n_0_0_26), .ZN(n_0_485));
   AOI222_X1 i_0_0_49 (.A1(n_0_422), .A2(n_0_0_39), .B1(n_0_438), .B2(n_0_0_38), 
      .C1(n_0_501), .C2(n_0_0_37), .ZN(n_0_0_26));
   INV_X1 i_0_0_50 (.A(n_0_0_27), .ZN(n_0_486));
   AOI222_X1 i_0_0_51 (.A1(n_0_423), .A2(n_0_0_39), .B1(n_0_439), .B2(n_0_0_38), 
      .C1(n_0_502), .C2(n_0_0_37), .ZN(n_0_0_27));
   INV_X1 i_0_0_52 (.A(n_0_0_28), .ZN(n_0_487));
   AOI222_X1 i_0_0_53 (.A1(n_0_424), .A2(n_0_0_39), .B1(n_0_440), .B2(n_0_0_38), 
      .C1(n_0_503), .C2(n_0_0_37), .ZN(n_0_0_28));
   INV_X1 i_0_0_54 (.A(n_0_0_29), .ZN(n_0_488));
   AOI222_X1 i_0_0_55 (.A1(n_0_425), .A2(n_0_0_39), .B1(n_0_441), .B2(n_0_0_38), 
      .C1(n_0_504), .C2(n_0_0_37), .ZN(n_0_0_29));
   INV_X1 i_0_0_56 (.A(n_0_0_30), .ZN(n_0_489));
   AOI222_X1 i_0_0_57 (.A1(n_0_426), .A2(n_0_0_39), .B1(n_0_442), .B2(n_0_0_38), 
      .C1(n_0_505), .C2(n_0_0_37), .ZN(n_0_0_30));
   INV_X1 i_0_0_58 (.A(n_0_0_31), .ZN(n_0_490));
   AOI222_X1 i_0_0_59 (.A1(n_0_427), .A2(n_0_0_39), .B1(n_0_443), .B2(n_0_0_38), 
      .C1(n_0_506), .C2(n_0_0_37), .ZN(n_0_0_31));
   INV_X1 i_0_0_60 (.A(n_0_0_32), .ZN(n_0_491));
   AOI222_X1 i_0_0_61 (.A1(n_0_428), .A2(n_0_0_39), .B1(n_0_444), .B2(n_0_0_38), 
      .C1(n_0_507), .C2(n_0_0_37), .ZN(n_0_0_32));
   INV_X1 i_0_0_62 (.A(n_0_0_33), .ZN(n_0_492));
   AOI222_X1 i_0_0_63 (.A1(n_0_429), .A2(n_0_0_39), .B1(n_0_445), .B2(n_0_0_38), 
      .C1(n_0_508), .C2(n_0_0_37), .ZN(n_0_0_33));
   INV_X1 i_0_0_64 (.A(n_0_0_34), .ZN(n_0_493));
   AOI221_X1 i_0_0_65 (.A(n_0_0_36), .B1(n_0_430), .B2(n_0_0_39), .C1(n_0_446), 
      .C2(n_0_0_38), .ZN(n_0_0_34));
   INV_X1 i_0_0_66 (.A(n_0_0_35), .ZN(n_0_494));
   AOI221_X1 i_0_0_67 (.A(n_0_0_36), .B1(n_0_431), .B2(n_0_0_39), .C1(n_0_447), 
      .C2(n_0_0_38), .ZN(n_0_0_35));
   AND2_X1 i_0_0_68 (.A1(n_0_509), .A2(n_0_0_37), .ZN(n_0_0_36));
   NOR2_X1 i_0_0_69 (.A1(n_0_0_39), .A2(n_0_0_38), .ZN(n_0_0_37));
   NOR2_X1 i_0_0_70 (.A1(multiplier[14]), .A2(n_0_0_340), .ZN(n_0_0_38));
   NOR2_X1 i_0_0_71 (.A1(n_0_0_341), .A2(multiplier[13]), .ZN(n_0_0_39));
   INV_X1 i_0_0_72 (.A(n_0_0_40), .ZN(product[13]));
   AOI222_X1 i_0_0_73 (.A1(n_0_400), .A2(n_0_0_59), .B1(n_0_384), .B2(n_0_0_58), 
      .C1(n_0_510), .C2(n_0_0_57), .ZN(n_0_0_40));
   INV_X1 i_0_0_74 (.A(n_0_0_41), .ZN(n_0_495));
   AOI222_X1 i_0_0_75 (.A1(n_0_401), .A2(n_0_0_59), .B1(n_0_385), .B2(n_0_0_58), 
      .C1(n_0_511), .C2(n_0_0_57), .ZN(n_0_0_41));
   INV_X1 i_0_0_76 (.A(n_0_0_42), .ZN(n_0_496));
   AOI222_X1 i_0_0_77 (.A1(n_0_402), .A2(n_0_0_59), .B1(n_0_386), .B2(n_0_0_58), 
      .C1(n_0_512), .C2(n_0_0_57), .ZN(n_0_0_42));
   INV_X1 i_0_0_78 (.A(n_0_0_43), .ZN(n_0_497));
   AOI222_X1 i_0_0_79 (.A1(n_0_403), .A2(n_0_0_59), .B1(n_0_387), .B2(n_0_0_58), 
      .C1(n_0_513), .C2(n_0_0_57), .ZN(n_0_0_43));
   INV_X1 i_0_0_80 (.A(n_0_0_44), .ZN(n_0_498));
   AOI222_X1 i_0_0_81 (.A1(n_0_404), .A2(n_0_0_59), .B1(n_0_388), .B2(n_0_0_58), 
      .C1(n_0_514), .C2(n_0_0_57), .ZN(n_0_0_44));
   INV_X1 i_0_0_82 (.A(n_0_0_45), .ZN(n_0_499));
   AOI222_X1 i_0_0_83 (.A1(n_0_405), .A2(n_0_0_59), .B1(n_0_389), .B2(n_0_0_58), 
      .C1(n_0_515), .C2(n_0_0_57), .ZN(n_0_0_45));
   INV_X1 i_0_0_84 (.A(n_0_0_46), .ZN(n_0_500));
   AOI222_X1 i_0_0_85 (.A1(n_0_406), .A2(n_0_0_59), .B1(n_0_390), .B2(n_0_0_58), 
      .C1(n_0_516), .C2(n_0_0_57), .ZN(n_0_0_46));
   INV_X1 i_0_0_86 (.A(n_0_0_47), .ZN(n_0_501));
   AOI222_X1 i_0_0_87 (.A1(n_0_407), .A2(n_0_0_59), .B1(n_0_391), .B2(n_0_0_58), 
      .C1(n_0_517), .C2(n_0_0_57), .ZN(n_0_0_47));
   INV_X1 i_0_0_88 (.A(n_0_0_48), .ZN(n_0_502));
   AOI222_X1 i_0_0_89 (.A1(n_0_408), .A2(n_0_0_59), .B1(n_0_392), .B2(n_0_0_58), 
      .C1(n_0_518), .C2(n_0_0_57), .ZN(n_0_0_48));
   INV_X1 i_0_0_90 (.A(n_0_0_49), .ZN(n_0_503));
   AOI222_X1 i_0_0_91 (.A1(n_0_409), .A2(n_0_0_59), .B1(n_0_393), .B2(n_0_0_58), 
      .C1(n_0_519), .C2(n_0_0_57), .ZN(n_0_0_49));
   INV_X1 i_0_0_92 (.A(n_0_0_50), .ZN(n_0_504));
   AOI222_X1 i_0_0_93 (.A1(n_0_410), .A2(n_0_0_59), .B1(n_0_394), .B2(n_0_0_58), 
      .C1(n_0_520), .C2(n_0_0_57), .ZN(n_0_0_50));
   INV_X1 i_0_0_94 (.A(n_0_0_51), .ZN(n_0_505));
   AOI222_X1 i_0_0_95 (.A1(n_0_411), .A2(n_0_0_59), .B1(n_0_395), .B2(n_0_0_58), 
      .C1(n_0_521), .C2(n_0_0_57), .ZN(n_0_0_51));
   INV_X1 i_0_0_96 (.A(n_0_0_52), .ZN(n_0_506));
   AOI222_X1 i_0_0_97 (.A1(n_0_412), .A2(n_0_0_59), .B1(n_0_396), .B2(n_0_0_58), 
      .C1(n_0_522), .C2(n_0_0_57), .ZN(n_0_0_52));
   INV_X1 i_0_0_98 (.A(n_0_0_53), .ZN(n_0_507));
   AOI222_X1 i_0_0_99 (.A1(n_0_413), .A2(n_0_0_59), .B1(n_0_397), .B2(n_0_0_58), 
      .C1(n_0_523), .C2(n_0_0_57), .ZN(n_0_0_53));
   INV_X1 i_0_0_100 (.A(n_0_0_54), .ZN(n_0_508));
   AOI221_X1 i_0_0_101 (.A(n_0_0_56), .B1(n_0_414), .B2(n_0_0_59), .C1(n_0_398), 
      .C2(n_0_0_58), .ZN(n_0_0_54));
   INV_X1 i_0_0_102 (.A(n_0_0_55), .ZN(n_0_509));
   AOI221_X1 i_0_0_103 (.A(n_0_0_56), .B1(n_0_415), .B2(n_0_0_59), .C1(n_0_399), 
      .C2(n_0_0_58), .ZN(n_0_0_55));
   AND2_X1 i_0_0_104 (.A1(n_0_524), .A2(n_0_0_57), .ZN(n_0_0_56));
   NOR2_X1 i_0_0_105 (.A1(n_0_0_59), .A2(n_0_0_58), .ZN(n_0_0_57));
   NOR2_X1 i_0_0_106 (.A1(n_0_0_340), .A2(multiplier[12]), .ZN(n_0_0_58));
   NOR2_X1 i_0_0_107 (.A1(multiplier[13]), .A2(n_0_0_339), .ZN(n_0_0_59));
   INV_X1 i_0_0_108 (.A(n_0_0_60), .ZN(product[12]));
   AOI222_X1 i_0_0_109 (.A1(n_0_368), .A2(n_0_0_79), .B1(n_0_352), .B2(n_0_0_78), 
      .C1(n_0_525), .C2(n_0_0_77), .ZN(n_0_0_60));
   INV_X1 i_0_0_110 (.A(n_0_0_61), .ZN(n_0_510));
   AOI222_X1 i_0_0_111 (.A1(n_0_369), .A2(n_0_0_79), .B1(n_0_353), .B2(n_0_0_78), 
      .C1(n_0_526), .C2(n_0_0_77), .ZN(n_0_0_61));
   INV_X1 i_0_0_112 (.A(n_0_0_62), .ZN(n_0_511));
   AOI222_X1 i_0_0_113 (.A1(n_0_370), .A2(n_0_0_79), .B1(n_0_354), .B2(n_0_0_78), 
      .C1(n_0_527), .C2(n_0_0_77), .ZN(n_0_0_62));
   INV_X1 i_0_0_114 (.A(n_0_0_63), .ZN(n_0_512));
   AOI222_X1 i_0_0_115 (.A1(n_0_371), .A2(n_0_0_79), .B1(n_0_355), .B2(n_0_0_78), 
      .C1(n_0_528), .C2(n_0_0_77), .ZN(n_0_0_63));
   INV_X1 i_0_0_116 (.A(n_0_0_64), .ZN(n_0_513));
   AOI222_X1 i_0_0_117 (.A1(n_0_372), .A2(n_0_0_79), .B1(n_0_356), .B2(n_0_0_78), 
      .C1(n_0_529), .C2(n_0_0_77), .ZN(n_0_0_64));
   INV_X1 i_0_0_118 (.A(n_0_0_65), .ZN(n_0_514));
   AOI222_X1 i_0_0_119 (.A1(n_0_373), .A2(n_0_0_79), .B1(n_0_357), .B2(n_0_0_78), 
      .C1(n_0_530), .C2(n_0_0_77), .ZN(n_0_0_65));
   INV_X1 i_0_0_120 (.A(n_0_0_66), .ZN(n_0_515));
   AOI222_X1 i_0_0_121 (.A1(n_0_374), .A2(n_0_0_79), .B1(n_0_358), .B2(n_0_0_78), 
      .C1(n_0_531), .C2(n_0_0_77), .ZN(n_0_0_66));
   INV_X1 i_0_0_122 (.A(n_0_0_67), .ZN(n_0_516));
   AOI222_X1 i_0_0_123 (.A1(n_0_375), .A2(n_0_0_79), .B1(n_0_359), .B2(n_0_0_78), 
      .C1(n_0_532), .C2(n_0_0_77), .ZN(n_0_0_67));
   INV_X1 i_0_0_124 (.A(n_0_0_68), .ZN(n_0_517));
   AOI222_X1 i_0_0_125 (.A1(n_0_376), .A2(n_0_0_79), .B1(n_0_360), .B2(n_0_0_78), 
      .C1(n_0_533), .C2(n_0_0_77), .ZN(n_0_0_68));
   INV_X1 i_0_0_126 (.A(n_0_0_69), .ZN(n_0_518));
   AOI222_X1 i_0_0_127 (.A1(n_0_377), .A2(n_0_0_79), .B1(n_0_361), .B2(n_0_0_78), 
      .C1(n_0_534), .C2(n_0_0_77), .ZN(n_0_0_69));
   INV_X1 i_0_0_128 (.A(n_0_0_70), .ZN(n_0_519));
   AOI222_X1 i_0_0_129 (.A1(n_0_378), .A2(n_0_0_79), .B1(n_0_362), .B2(n_0_0_78), 
      .C1(n_0_535), .C2(n_0_0_77), .ZN(n_0_0_70));
   INV_X1 i_0_0_130 (.A(n_0_0_71), .ZN(n_0_520));
   AOI222_X1 i_0_0_131 (.A1(n_0_379), .A2(n_0_0_79), .B1(n_0_363), .B2(n_0_0_78), 
      .C1(n_0_536), .C2(n_0_0_77), .ZN(n_0_0_71));
   INV_X1 i_0_0_132 (.A(n_0_0_72), .ZN(n_0_521));
   AOI222_X1 i_0_0_133 (.A1(n_0_380), .A2(n_0_0_79), .B1(n_0_364), .B2(n_0_0_78), 
      .C1(n_0_537), .C2(n_0_0_77), .ZN(n_0_0_72));
   INV_X1 i_0_0_134 (.A(n_0_0_73), .ZN(n_0_522));
   AOI222_X1 i_0_0_135 (.A1(n_0_381), .A2(n_0_0_79), .B1(n_0_365), .B2(n_0_0_78), 
      .C1(n_0_538), .C2(n_0_0_77), .ZN(n_0_0_73));
   INV_X1 i_0_0_136 (.A(n_0_0_74), .ZN(n_0_523));
   AOI221_X1 i_0_0_137 (.A(n_0_0_76), .B1(n_0_382), .B2(n_0_0_79), .C1(n_0_366), 
      .C2(n_0_0_78), .ZN(n_0_0_74));
   INV_X1 i_0_0_138 (.A(n_0_0_75), .ZN(n_0_524));
   AOI221_X1 i_0_0_139 (.A(n_0_0_76), .B1(n_0_383), .B2(n_0_0_79), .C1(n_0_367), 
      .C2(n_0_0_78), .ZN(n_0_0_75));
   AND2_X1 i_0_0_140 (.A1(n_0_539), .A2(n_0_0_77), .ZN(n_0_0_76));
   NOR2_X1 i_0_0_141 (.A1(n_0_0_79), .A2(n_0_0_78), .ZN(n_0_0_77));
   NOR2_X1 i_0_0_142 (.A1(n_0_0_339), .A2(multiplier[11]), .ZN(n_0_0_78));
   NOR2_X1 i_0_0_143 (.A1(multiplier[12]), .A2(n_0_0_338), .ZN(n_0_0_79));
   INV_X1 i_0_0_144 (.A(n_0_0_80), .ZN(product[11]));
   AOI222_X1 i_0_0_145 (.A1(n_0_320), .A2(n_0_0_98), .B1(n_0_336), .B2(n_0_0_99), 
      .C1(n_0_540), .C2(n_0_0_97), .ZN(n_0_0_80));
   INV_X1 i_0_0_146 (.A(n_0_0_81), .ZN(n_0_525));
   AOI222_X1 i_0_0_147 (.A1(n_0_321), .A2(n_0_0_98), .B1(n_0_337), .B2(n_0_0_99), 
      .C1(n_0_541), .C2(n_0_0_97), .ZN(n_0_0_81));
   INV_X1 i_0_0_148 (.A(n_0_0_82), .ZN(n_0_526));
   AOI222_X1 i_0_0_149 (.A1(n_0_338), .A2(n_0_0_99), .B1(n_0_322), .B2(n_0_0_98), 
      .C1(n_0_542), .C2(n_0_0_97), .ZN(n_0_0_82));
   INV_X1 i_0_0_150 (.A(n_0_0_83), .ZN(n_0_527));
   AOI222_X1 i_0_0_151 (.A1(n_0_339), .A2(n_0_0_99), .B1(n_0_323), .B2(n_0_0_98), 
      .C1(n_0_543), .C2(n_0_0_97), .ZN(n_0_0_83));
   INV_X1 i_0_0_152 (.A(n_0_0_84), .ZN(n_0_528));
   AOI222_X1 i_0_0_153 (.A1(n_0_340), .A2(n_0_0_99), .B1(n_0_324), .B2(n_0_0_98), 
      .C1(n_0_544), .C2(n_0_0_97), .ZN(n_0_0_84));
   INV_X1 i_0_0_154 (.A(n_0_0_85), .ZN(n_0_529));
   AOI222_X1 i_0_0_155 (.A1(n_0_341), .A2(n_0_0_99), .B1(n_0_325), .B2(n_0_0_98), 
      .C1(n_0_545), .C2(n_0_0_97), .ZN(n_0_0_85));
   INV_X1 i_0_0_156 (.A(n_0_0_86), .ZN(n_0_530));
   AOI222_X1 i_0_0_157 (.A1(n_0_342), .A2(n_0_0_99), .B1(n_0_326), .B2(n_0_0_98), 
      .C1(n_0_546), .C2(n_0_0_97), .ZN(n_0_0_86));
   INV_X1 i_0_0_158 (.A(n_0_0_87), .ZN(n_0_531));
   AOI222_X1 i_0_0_159 (.A1(n_0_343), .A2(n_0_0_99), .B1(n_0_327), .B2(n_0_0_98), 
      .C1(n_0_547), .C2(n_0_0_97), .ZN(n_0_0_87));
   INV_X1 i_0_0_160 (.A(n_0_0_88), .ZN(n_0_532));
   AOI222_X1 i_0_0_161 (.A1(n_0_344), .A2(n_0_0_99), .B1(n_0_328), .B2(n_0_0_98), 
      .C1(n_0_548), .C2(n_0_0_97), .ZN(n_0_0_88));
   INV_X1 i_0_0_162 (.A(n_0_0_89), .ZN(n_0_533));
   AOI222_X1 i_0_0_163 (.A1(n_0_345), .A2(n_0_0_99), .B1(n_0_329), .B2(n_0_0_98), 
      .C1(n_0_549), .C2(n_0_0_97), .ZN(n_0_0_89));
   INV_X1 i_0_0_164 (.A(n_0_0_90), .ZN(n_0_534));
   AOI222_X1 i_0_0_165 (.A1(n_0_346), .A2(n_0_0_99), .B1(n_0_330), .B2(n_0_0_98), 
      .C1(n_0_550), .C2(n_0_0_97), .ZN(n_0_0_90));
   INV_X1 i_0_0_166 (.A(n_0_0_91), .ZN(n_0_535));
   AOI222_X1 i_0_0_167 (.A1(n_0_347), .A2(n_0_0_99), .B1(n_0_331), .B2(n_0_0_98), 
      .C1(n_0_551), .C2(n_0_0_97), .ZN(n_0_0_91));
   INV_X1 i_0_0_168 (.A(n_0_0_92), .ZN(n_0_536));
   AOI222_X1 i_0_0_169 (.A1(n_0_348), .A2(n_0_0_99), .B1(n_0_332), .B2(n_0_0_98), 
      .C1(n_0_552), .C2(n_0_0_97), .ZN(n_0_0_92));
   INV_X1 i_0_0_170 (.A(n_0_0_93), .ZN(n_0_537));
   AOI222_X1 i_0_0_171 (.A1(n_0_349), .A2(n_0_0_99), .B1(n_0_333), .B2(n_0_0_98), 
      .C1(n_0_553), .C2(n_0_0_97), .ZN(n_0_0_93));
   INV_X1 i_0_0_172 (.A(n_0_0_94), .ZN(n_0_538));
   AOI221_X1 i_0_0_173 (.A(n_0_0_96), .B1(n_0_350), .B2(n_0_0_99), .C1(n_0_334), 
      .C2(n_0_0_98), .ZN(n_0_0_94));
   INV_X1 i_0_0_174 (.A(n_0_0_95), .ZN(n_0_539));
   AOI221_X1 i_0_0_175 (.A(n_0_0_96), .B1(n_0_351), .B2(n_0_0_99), .C1(n_0_335), 
      .C2(n_0_0_98), .ZN(n_0_0_95));
   AND2_X1 i_0_0_176 (.A1(n_0_554), .A2(n_0_0_97), .ZN(n_0_0_96));
   NOR2_X1 i_0_0_177 (.A1(n_0_0_99), .A2(n_0_0_98), .ZN(n_0_0_97));
   NOR2_X1 i_0_0_178 (.A1(n_0_0_338), .A2(multiplier[10]), .ZN(n_0_0_98));
   NOR2_X1 i_0_0_179 (.A1(multiplier[11]), .A2(n_0_0_337), .ZN(n_0_0_99));
   INV_X1 i_0_0_180 (.A(n_0_0_100), .ZN(product[10]));
   AOI222_X1 i_0_0_181 (.A1(n_0_288), .A2(n_0_0_118), .B1(n_0_304), .B2(
      n_0_0_119), .C1(n_0_555), .C2(n_0_0_117), .ZN(n_0_0_100));
   INV_X1 i_0_0_182 (.A(n_0_0_101), .ZN(n_0_540));
   AOI222_X1 i_0_0_183 (.A1(n_0_289), .A2(n_0_0_118), .B1(n_0_305), .B2(
      n_0_0_119), .C1(n_0_556), .C2(n_0_0_117), .ZN(n_0_0_101));
   INV_X1 i_0_0_184 (.A(n_0_0_102), .ZN(n_0_541));
   AOI222_X1 i_0_0_185 (.A1(n_0_290), .A2(n_0_0_118), .B1(n_0_306), .B2(
      n_0_0_119), .C1(n_0_557), .C2(n_0_0_117), .ZN(n_0_0_102));
   INV_X1 i_0_0_186 (.A(n_0_0_103), .ZN(n_0_542));
   AOI222_X1 i_0_0_187 (.A1(n_0_307), .A2(n_0_0_119), .B1(n_0_291), .B2(
      n_0_0_118), .C1(n_0_558), .C2(n_0_0_117), .ZN(n_0_0_103));
   INV_X1 i_0_0_188 (.A(n_0_0_104), .ZN(n_0_543));
   AOI222_X1 i_0_0_189 (.A1(n_0_308), .A2(n_0_0_119), .B1(n_0_292), .B2(
      n_0_0_118), .C1(n_0_559), .C2(n_0_0_117), .ZN(n_0_0_104));
   INV_X1 i_0_0_190 (.A(n_0_0_105), .ZN(n_0_544));
   AOI222_X1 i_0_0_191 (.A1(n_0_309), .A2(n_0_0_119), .B1(n_0_293), .B2(
      n_0_0_118), .C1(n_0_560), .C2(n_0_0_117), .ZN(n_0_0_105));
   INV_X1 i_0_0_192 (.A(n_0_0_106), .ZN(n_0_545));
   AOI222_X1 i_0_0_193 (.A1(n_0_310), .A2(n_0_0_119), .B1(n_0_294), .B2(
      n_0_0_118), .C1(n_0_561), .C2(n_0_0_117), .ZN(n_0_0_106));
   INV_X1 i_0_0_194 (.A(n_0_0_107), .ZN(n_0_546));
   AOI222_X1 i_0_0_195 (.A1(n_0_311), .A2(n_0_0_119), .B1(n_0_295), .B2(
      n_0_0_118), .C1(n_0_562), .C2(n_0_0_117), .ZN(n_0_0_107));
   INV_X1 i_0_0_196 (.A(n_0_0_108), .ZN(n_0_547));
   AOI222_X1 i_0_0_197 (.A1(n_0_312), .A2(n_0_0_119), .B1(n_0_296), .B2(
      n_0_0_118), .C1(n_0_563), .C2(n_0_0_117), .ZN(n_0_0_108));
   INV_X1 i_0_0_198 (.A(n_0_0_109), .ZN(n_0_548));
   AOI222_X1 i_0_0_199 (.A1(n_0_313), .A2(n_0_0_119), .B1(n_0_297), .B2(
      n_0_0_118), .C1(n_0_564), .C2(n_0_0_117), .ZN(n_0_0_109));
   INV_X1 i_0_0_200 (.A(n_0_0_110), .ZN(n_0_549));
   AOI222_X1 i_0_0_201 (.A1(n_0_314), .A2(n_0_0_119), .B1(n_0_298), .B2(
      n_0_0_118), .C1(n_0_565), .C2(n_0_0_117), .ZN(n_0_0_110));
   INV_X1 i_0_0_202 (.A(n_0_0_111), .ZN(n_0_550));
   AOI222_X1 i_0_0_203 (.A1(n_0_315), .A2(n_0_0_119), .B1(n_0_299), .B2(
      n_0_0_118), .C1(n_0_566), .C2(n_0_0_117), .ZN(n_0_0_111));
   INV_X1 i_0_0_204 (.A(n_0_0_112), .ZN(n_0_551));
   AOI222_X1 i_0_0_205 (.A1(n_0_316), .A2(n_0_0_119), .B1(n_0_300), .B2(
      n_0_0_118), .C1(n_0_567), .C2(n_0_0_117), .ZN(n_0_0_112));
   INV_X1 i_0_0_206 (.A(n_0_0_113), .ZN(n_0_552));
   AOI222_X1 i_0_0_207 (.A1(n_0_317), .A2(n_0_0_119), .B1(n_0_301), .B2(
      n_0_0_118), .C1(n_0_568), .C2(n_0_0_117), .ZN(n_0_0_113));
   INV_X1 i_0_0_208 (.A(n_0_0_114), .ZN(n_0_553));
   AOI221_X1 i_0_0_209 (.A(n_0_0_116), .B1(n_0_318), .B2(n_0_0_119), .C1(n_0_302), 
      .C2(n_0_0_118), .ZN(n_0_0_114));
   INV_X1 i_0_0_210 (.A(n_0_0_115), .ZN(n_0_554));
   AOI221_X1 i_0_0_211 (.A(n_0_0_116), .B1(n_0_319), .B2(n_0_0_119), .C1(n_0_303), 
      .C2(n_0_0_118), .ZN(n_0_0_115));
   AND2_X1 i_0_0_212 (.A1(n_0_569), .A2(n_0_0_117), .ZN(n_0_0_116));
   NOR2_X1 i_0_0_213 (.A1(n_0_0_119), .A2(n_0_0_118), .ZN(n_0_0_117));
   NOR2_X1 i_0_0_214 (.A1(n_0_0_337), .A2(multiplier[9]), .ZN(n_0_0_118));
   NOR2_X1 i_0_0_215 (.A1(multiplier[10]), .A2(n_0_0_336), .ZN(n_0_0_119));
   INV_X1 i_0_0_216 (.A(n_0_0_120), .ZN(product[9]));
   AOI222_X1 i_0_0_217 (.A1(n_0_256), .A2(n_0_0_138), .B1(n_0_272), .B2(
      n_0_0_139), .C1(n_0_570), .C2(n_0_0_137), .ZN(n_0_0_120));
   INV_X1 i_0_0_218 (.A(n_0_0_121), .ZN(n_0_555));
   AOI222_X1 i_0_0_219 (.A1(n_0_257), .A2(n_0_0_138), .B1(n_0_273), .B2(
      n_0_0_139), .C1(n_0_571), .C2(n_0_0_137), .ZN(n_0_0_121));
   INV_X1 i_0_0_220 (.A(n_0_0_122), .ZN(n_0_556));
   AOI222_X1 i_0_0_221 (.A1(n_0_258), .A2(n_0_0_138), .B1(n_0_274), .B2(
      n_0_0_139), .C1(n_0_572), .C2(n_0_0_137), .ZN(n_0_0_122));
   INV_X1 i_0_0_222 (.A(n_0_0_123), .ZN(n_0_557));
   AOI222_X1 i_0_0_223 (.A1(n_0_259), .A2(n_0_0_138), .B1(n_0_275), .B2(
      n_0_0_139), .C1(n_0_573), .C2(n_0_0_137), .ZN(n_0_0_123));
   INV_X1 i_0_0_224 (.A(n_0_0_124), .ZN(n_0_558));
   AOI222_X1 i_0_0_225 (.A1(n_0_276), .A2(n_0_0_139), .B1(n_0_260), .B2(
      n_0_0_138), .C1(n_0_574), .C2(n_0_0_137), .ZN(n_0_0_124));
   INV_X1 i_0_0_226 (.A(n_0_0_125), .ZN(n_0_559));
   AOI222_X1 i_0_0_227 (.A1(n_0_277), .A2(n_0_0_139), .B1(n_0_261), .B2(
      n_0_0_138), .C1(n_0_575), .C2(n_0_0_137), .ZN(n_0_0_125));
   INV_X1 i_0_0_228 (.A(n_0_0_126), .ZN(n_0_560));
   AOI222_X1 i_0_0_229 (.A1(n_0_278), .A2(n_0_0_139), .B1(n_0_262), .B2(
      n_0_0_138), .C1(n_0_576), .C2(n_0_0_137), .ZN(n_0_0_126));
   INV_X1 i_0_0_230 (.A(n_0_0_127), .ZN(n_0_561));
   AOI222_X1 i_0_0_231 (.A1(n_0_279), .A2(n_0_0_139), .B1(n_0_263), .B2(
      n_0_0_138), .C1(n_0_577), .C2(n_0_0_137), .ZN(n_0_0_127));
   INV_X1 i_0_0_232 (.A(n_0_0_128), .ZN(n_0_562));
   AOI222_X1 i_0_0_233 (.A1(n_0_280), .A2(n_0_0_139), .B1(n_0_264), .B2(
      n_0_0_138), .C1(n_0_578), .C2(n_0_0_137), .ZN(n_0_0_128));
   INV_X1 i_0_0_234 (.A(n_0_0_129), .ZN(n_0_563));
   AOI222_X1 i_0_0_235 (.A1(n_0_281), .A2(n_0_0_139), .B1(n_0_265), .B2(
      n_0_0_138), .C1(n_0_579), .C2(n_0_0_137), .ZN(n_0_0_129));
   INV_X1 i_0_0_236 (.A(n_0_0_130), .ZN(n_0_564));
   AOI222_X1 i_0_0_237 (.A1(n_0_282), .A2(n_0_0_139), .B1(n_0_266), .B2(
      n_0_0_138), .C1(n_0_580), .C2(n_0_0_137), .ZN(n_0_0_130));
   INV_X1 i_0_0_238 (.A(n_0_0_131), .ZN(n_0_565));
   AOI222_X1 i_0_0_239 (.A1(n_0_283), .A2(n_0_0_139), .B1(n_0_267), .B2(
      n_0_0_138), .C1(n_0_581), .C2(n_0_0_137), .ZN(n_0_0_131));
   INV_X1 i_0_0_240 (.A(n_0_0_132), .ZN(n_0_566));
   AOI222_X1 i_0_0_241 (.A1(n_0_284), .A2(n_0_0_139), .B1(n_0_268), .B2(
      n_0_0_138), .C1(n_0_582), .C2(n_0_0_137), .ZN(n_0_0_132));
   INV_X1 i_0_0_242 (.A(n_0_0_133), .ZN(n_0_567));
   AOI222_X1 i_0_0_243 (.A1(n_0_285), .A2(n_0_0_139), .B1(n_0_269), .B2(
      n_0_0_138), .C1(n_0_583), .C2(n_0_0_137), .ZN(n_0_0_133));
   INV_X1 i_0_0_244 (.A(n_0_0_134), .ZN(n_0_568));
   AOI221_X1 i_0_0_245 (.A(n_0_0_136), .B1(n_0_286), .B2(n_0_0_139), .C1(n_0_270), 
      .C2(n_0_0_138), .ZN(n_0_0_134));
   INV_X1 i_0_0_246 (.A(n_0_0_135), .ZN(n_0_569));
   AOI221_X1 i_0_0_247 (.A(n_0_0_136), .B1(n_0_287), .B2(n_0_0_139), .C1(n_0_271), 
      .C2(n_0_0_138), .ZN(n_0_0_135));
   AND2_X1 i_0_0_248 (.A1(n_0_584), .A2(n_0_0_137), .ZN(n_0_0_136));
   NOR2_X1 i_0_0_249 (.A1(n_0_0_139), .A2(n_0_0_138), .ZN(n_0_0_137));
   NOR2_X1 i_0_0_250 (.A1(n_0_0_336), .A2(multiplier[8]), .ZN(n_0_0_138));
   NOR2_X1 i_0_0_251 (.A1(multiplier[9]), .A2(n_0_0_335), .ZN(n_0_0_139));
   INV_X1 i_0_0_252 (.A(n_0_0_140), .ZN(product[8]));
   AOI222_X1 i_0_0_253 (.A1(n_0_224), .A2(n_0_0_158), .B1(n_0_240), .B2(
      n_0_0_159), .C1(n_0_585), .C2(n_0_0_157), .ZN(n_0_0_140));
   INV_X1 i_0_0_254 (.A(n_0_0_141), .ZN(n_0_570));
   AOI222_X1 i_0_0_255 (.A1(n_0_225), .A2(n_0_0_158), .B1(n_0_241), .B2(
      n_0_0_159), .C1(n_0_586), .C2(n_0_0_157), .ZN(n_0_0_141));
   INV_X1 i_0_0_256 (.A(n_0_0_142), .ZN(n_0_571));
   AOI222_X1 i_0_0_257 (.A1(n_0_226), .A2(n_0_0_158), .B1(n_0_242), .B2(
      n_0_0_159), .C1(n_0_587), .C2(n_0_0_157), .ZN(n_0_0_142));
   INV_X1 i_0_0_258 (.A(n_0_0_143), .ZN(n_0_572));
   AOI222_X1 i_0_0_259 (.A1(n_0_227), .A2(n_0_0_158), .B1(n_0_243), .B2(
      n_0_0_159), .C1(n_0_588), .C2(n_0_0_157), .ZN(n_0_0_143));
   INV_X1 i_0_0_260 (.A(n_0_0_144), .ZN(n_0_573));
   AOI222_X1 i_0_0_261 (.A1(n_0_228), .A2(n_0_0_158), .B1(n_0_244), .B2(
      n_0_0_159), .C1(n_0_589), .C2(n_0_0_157), .ZN(n_0_0_144));
   INV_X1 i_0_0_262 (.A(n_0_0_145), .ZN(n_0_574));
   AOI222_X1 i_0_0_263 (.A1(n_0_229), .A2(n_0_0_158), .B1(n_0_245), .B2(
      n_0_0_159), .C1(n_0_590), .C2(n_0_0_157), .ZN(n_0_0_145));
   INV_X1 i_0_0_264 (.A(n_0_0_146), .ZN(n_0_575));
   AOI222_X1 i_0_0_265 (.A1(n_0_246), .A2(n_0_0_159), .B1(n_0_230), .B2(
      n_0_0_158), .C1(n_0_591), .C2(n_0_0_157), .ZN(n_0_0_146));
   INV_X1 i_0_0_266 (.A(n_0_0_147), .ZN(n_0_576));
   AOI222_X1 i_0_0_267 (.A1(n_0_247), .A2(n_0_0_159), .B1(n_0_231), .B2(
      n_0_0_158), .C1(n_0_592), .C2(n_0_0_157), .ZN(n_0_0_147));
   INV_X1 i_0_0_268 (.A(n_0_0_148), .ZN(n_0_577));
   AOI222_X1 i_0_0_269 (.A1(n_0_248), .A2(n_0_0_159), .B1(n_0_232), .B2(
      n_0_0_158), .C1(n_0_593), .C2(n_0_0_157), .ZN(n_0_0_148));
   INV_X1 i_0_0_270 (.A(n_0_0_149), .ZN(n_0_578));
   AOI222_X1 i_0_0_271 (.A1(n_0_249), .A2(n_0_0_159), .B1(n_0_233), .B2(
      n_0_0_158), .C1(n_0_594), .C2(n_0_0_157), .ZN(n_0_0_149));
   INV_X1 i_0_0_272 (.A(n_0_0_150), .ZN(n_0_579));
   AOI222_X1 i_0_0_273 (.A1(n_0_250), .A2(n_0_0_159), .B1(n_0_234), .B2(
      n_0_0_158), .C1(n_0_595), .C2(n_0_0_157), .ZN(n_0_0_150));
   INV_X1 i_0_0_274 (.A(n_0_0_151), .ZN(n_0_580));
   AOI222_X1 i_0_0_275 (.A1(n_0_251), .A2(n_0_0_159), .B1(n_0_235), .B2(
      n_0_0_158), .C1(n_0_596), .C2(n_0_0_157), .ZN(n_0_0_151));
   INV_X1 i_0_0_276 (.A(n_0_0_152), .ZN(n_0_581));
   AOI222_X1 i_0_0_277 (.A1(n_0_252), .A2(n_0_0_159), .B1(n_0_236), .B2(
      n_0_0_158), .C1(n_0_597), .C2(n_0_0_157), .ZN(n_0_0_152));
   INV_X1 i_0_0_278 (.A(n_0_0_153), .ZN(n_0_582));
   AOI222_X1 i_0_0_279 (.A1(n_0_253), .A2(n_0_0_159), .B1(n_0_237), .B2(
      n_0_0_158), .C1(n_0_598), .C2(n_0_0_157), .ZN(n_0_0_153));
   INV_X1 i_0_0_280 (.A(n_0_0_154), .ZN(n_0_583));
   AOI221_X1 i_0_0_281 (.A(n_0_0_156), .B1(n_0_254), .B2(n_0_0_159), .C1(n_0_238), 
      .C2(n_0_0_158), .ZN(n_0_0_154));
   INV_X1 i_0_0_282 (.A(n_0_0_155), .ZN(n_0_584));
   AOI221_X1 i_0_0_283 (.A(n_0_0_156), .B1(n_0_255), .B2(n_0_0_159), .C1(n_0_239), 
      .C2(n_0_0_158), .ZN(n_0_0_155));
   AND2_X1 i_0_0_284 (.A1(n_0_599), .A2(n_0_0_157), .ZN(n_0_0_156));
   NOR2_X1 i_0_0_285 (.A1(n_0_0_159), .A2(n_0_0_158), .ZN(n_0_0_157));
   NOR2_X1 i_0_0_286 (.A1(n_0_0_335), .A2(multiplier[7]), .ZN(n_0_0_158));
   NOR2_X1 i_0_0_287 (.A1(multiplier[8]), .A2(n_0_0_334), .ZN(n_0_0_159));
   INV_X1 i_0_0_288 (.A(n_0_0_160), .ZN(product[7]));
   AOI222_X1 i_0_0_289 (.A1(n_0_192), .A2(n_0_0_178), .B1(n_0_208), .B2(
      n_0_0_179), .C1(n_0_600), .C2(n_0_0_177), .ZN(n_0_0_160));
   INV_X1 i_0_0_290 (.A(n_0_0_161), .ZN(n_0_585));
   AOI222_X1 i_0_0_291 (.A1(n_0_193), .A2(n_0_0_178), .B1(n_0_209), .B2(
      n_0_0_179), .C1(n_0_601), .C2(n_0_0_177), .ZN(n_0_0_161));
   INV_X1 i_0_0_292 (.A(n_0_0_162), .ZN(n_0_586));
   AOI222_X1 i_0_0_293 (.A1(n_0_194), .A2(n_0_0_178), .B1(n_0_210), .B2(
      n_0_0_179), .C1(n_0_602), .C2(n_0_0_177), .ZN(n_0_0_162));
   INV_X1 i_0_0_294 (.A(n_0_0_163), .ZN(n_0_587));
   AOI222_X1 i_0_0_295 (.A1(n_0_195), .A2(n_0_0_178), .B1(n_0_211), .B2(
      n_0_0_179), .C1(n_0_603), .C2(n_0_0_177), .ZN(n_0_0_163));
   INV_X1 i_0_0_296 (.A(n_0_0_164), .ZN(n_0_588));
   AOI222_X1 i_0_0_297 (.A1(n_0_196), .A2(n_0_0_178), .B1(n_0_212), .B2(
      n_0_0_179), .C1(n_0_604), .C2(n_0_0_177), .ZN(n_0_0_164));
   INV_X1 i_0_0_298 (.A(n_0_0_165), .ZN(n_0_589));
   AOI222_X1 i_0_0_299 (.A1(n_0_197), .A2(n_0_0_178), .B1(n_0_213), .B2(
      n_0_0_179), .C1(n_0_605), .C2(n_0_0_177), .ZN(n_0_0_165));
   INV_X1 i_0_0_300 (.A(n_0_0_166), .ZN(n_0_590));
   AOI222_X1 i_0_0_301 (.A1(n_0_198), .A2(n_0_0_178), .B1(n_0_214), .B2(
      n_0_0_179), .C1(n_0_606), .C2(n_0_0_177), .ZN(n_0_0_166));
   INV_X1 i_0_0_302 (.A(n_0_0_167), .ZN(n_0_591));
   AOI222_X1 i_0_0_303 (.A1(n_0_215), .A2(n_0_0_179), .B1(n_0_199), .B2(
      n_0_0_178), .C1(n_0_607), .C2(n_0_0_177), .ZN(n_0_0_167));
   INV_X1 i_0_0_304 (.A(n_0_0_168), .ZN(n_0_592));
   AOI222_X1 i_0_0_305 (.A1(n_0_216), .A2(n_0_0_179), .B1(n_0_200), .B2(
      n_0_0_178), .C1(n_0_608), .C2(n_0_0_177), .ZN(n_0_0_168));
   INV_X1 i_0_0_306 (.A(n_0_0_169), .ZN(n_0_593));
   AOI222_X1 i_0_0_307 (.A1(n_0_217), .A2(n_0_0_179), .B1(n_0_201), .B2(
      n_0_0_178), .C1(n_0_609), .C2(n_0_0_177), .ZN(n_0_0_169));
   INV_X1 i_0_0_308 (.A(n_0_0_170), .ZN(n_0_594));
   AOI222_X1 i_0_0_309 (.A1(n_0_218), .A2(n_0_0_179), .B1(n_0_202), .B2(
      n_0_0_178), .C1(n_0_610), .C2(n_0_0_177), .ZN(n_0_0_170));
   INV_X1 i_0_0_310 (.A(n_0_0_171), .ZN(n_0_595));
   AOI222_X1 i_0_0_311 (.A1(n_0_219), .A2(n_0_0_179), .B1(n_0_203), .B2(
      n_0_0_178), .C1(n_0_611), .C2(n_0_0_177), .ZN(n_0_0_171));
   INV_X1 i_0_0_312 (.A(n_0_0_172), .ZN(n_0_596));
   AOI222_X1 i_0_0_313 (.A1(n_0_220), .A2(n_0_0_179), .B1(n_0_204), .B2(
      n_0_0_178), .C1(n_0_612), .C2(n_0_0_177), .ZN(n_0_0_172));
   INV_X1 i_0_0_314 (.A(n_0_0_173), .ZN(n_0_597));
   AOI222_X1 i_0_0_315 (.A1(n_0_221), .A2(n_0_0_179), .B1(n_0_205), .B2(
      n_0_0_178), .C1(n_0_613), .C2(n_0_0_177), .ZN(n_0_0_173));
   INV_X1 i_0_0_316 (.A(n_0_0_174), .ZN(n_0_598));
   AOI221_X1 i_0_0_317 (.A(n_0_0_176), .B1(n_0_222), .B2(n_0_0_179), .C1(n_0_206), 
      .C2(n_0_0_178), .ZN(n_0_0_174));
   INV_X1 i_0_0_318 (.A(n_0_0_175), .ZN(n_0_599));
   AOI221_X1 i_0_0_319 (.A(n_0_0_176), .B1(n_0_223), .B2(n_0_0_179), .C1(n_0_207), 
      .C2(n_0_0_178), .ZN(n_0_0_175));
   AND2_X1 i_0_0_320 (.A1(n_0_614), .A2(n_0_0_177), .ZN(n_0_0_176));
   NOR2_X1 i_0_0_321 (.A1(n_0_0_179), .A2(n_0_0_178), .ZN(n_0_0_177));
   NOR2_X1 i_0_0_322 (.A1(n_0_0_334), .A2(multiplier[6]), .ZN(n_0_0_178));
   NOR2_X1 i_0_0_323 (.A1(multiplier[7]), .A2(n_0_0_333), .ZN(n_0_0_179));
   INV_X1 i_0_0_324 (.A(n_0_0_180), .ZN(product[6]));
   AOI222_X1 i_0_0_325 (.A1(n_0_160), .A2(n_0_0_198), .B1(n_0_176), .B2(
      n_0_0_199), .C1(n_0_615), .C2(n_0_0_197), .ZN(n_0_0_180));
   INV_X1 i_0_0_326 (.A(n_0_0_181), .ZN(n_0_600));
   AOI222_X1 i_0_0_327 (.A1(n_0_161), .A2(n_0_0_198), .B1(n_0_177), .B2(
      n_0_0_199), .C1(n_0_616), .C2(n_0_0_197), .ZN(n_0_0_181));
   INV_X1 i_0_0_328 (.A(n_0_0_182), .ZN(n_0_601));
   AOI222_X1 i_0_0_329 (.A1(n_0_162), .A2(n_0_0_198), .B1(n_0_178), .B2(
      n_0_0_199), .C1(n_0_617), .C2(n_0_0_197), .ZN(n_0_0_182));
   INV_X1 i_0_0_330 (.A(n_0_0_183), .ZN(n_0_602));
   AOI222_X1 i_0_0_331 (.A1(n_0_163), .A2(n_0_0_198), .B1(n_0_179), .B2(
      n_0_0_199), .C1(n_0_618), .C2(n_0_0_197), .ZN(n_0_0_183));
   INV_X1 i_0_0_332 (.A(n_0_0_184), .ZN(n_0_603));
   AOI222_X1 i_0_0_333 (.A1(n_0_164), .A2(n_0_0_198), .B1(n_0_180), .B2(
      n_0_0_199), .C1(n_0_619), .C2(n_0_0_197), .ZN(n_0_0_184));
   INV_X1 i_0_0_334 (.A(n_0_0_185), .ZN(n_0_604));
   AOI222_X1 i_0_0_335 (.A1(n_0_165), .A2(n_0_0_198), .B1(n_0_181), .B2(
      n_0_0_199), .C1(n_0_620), .C2(n_0_0_197), .ZN(n_0_0_185));
   INV_X1 i_0_0_336 (.A(n_0_0_186), .ZN(n_0_605));
   AOI222_X1 i_0_0_337 (.A1(n_0_166), .A2(n_0_0_198), .B1(n_0_182), .B2(
      n_0_0_199), .C1(n_0_621), .C2(n_0_0_197), .ZN(n_0_0_186));
   INV_X1 i_0_0_338 (.A(n_0_0_187), .ZN(n_0_606));
   AOI222_X1 i_0_0_339 (.A1(n_0_167), .A2(n_0_0_198), .B1(n_0_183), .B2(
      n_0_0_199), .C1(n_0_622), .C2(n_0_0_197), .ZN(n_0_0_187));
   INV_X1 i_0_0_340 (.A(n_0_0_188), .ZN(n_0_607));
   AOI222_X1 i_0_0_341 (.A1(n_0_184), .A2(n_0_0_199), .B1(n_0_168), .B2(
      n_0_0_198), .C1(n_0_623), .C2(n_0_0_197), .ZN(n_0_0_188));
   INV_X1 i_0_0_342 (.A(n_0_0_189), .ZN(n_0_608));
   AOI222_X1 i_0_0_343 (.A1(n_0_185), .A2(n_0_0_199), .B1(n_0_169), .B2(
      n_0_0_198), .C1(n_0_624), .C2(n_0_0_197), .ZN(n_0_0_189));
   INV_X1 i_0_0_344 (.A(n_0_0_190), .ZN(n_0_609));
   AOI222_X1 i_0_0_345 (.A1(n_0_186), .A2(n_0_0_199), .B1(n_0_170), .B2(
      n_0_0_198), .C1(n_0_625), .C2(n_0_0_197), .ZN(n_0_0_190));
   INV_X1 i_0_0_346 (.A(n_0_0_191), .ZN(n_0_610));
   AOI222_X1 i_0_0_347 (.A1(n_0_187), .A2(n_0_0_199), .B1(n_0_171), .B2(
      n_0_0_198), .C1(n_0_626), .C2(n_0_0_197), .ZN(n_0_0_191));
   INV_X1 i_0_0_348 (.A(n_0_0_192), .ZN(n_0_611));
   AOI222_X1 i_0_0_349 (.A1(n_0_188), .A2(n_0_0_199), .B1(n_0_172), .B2(
      n_0_0_198), .C1(n_0_627), .C2(n_0_0_197), .ZN(n_0_0_192));
   INV_X1 i_0_0_350 (.A(n_0_0_193), .ZN(n_0_612));
   AOI222_X1 i_0_0_351 (.A1(n_0_189), .A2(n_0_0_199), .B1(n_0_173), .B2(
      n_0_0_198), .C1(n_0_628), .C2(n_0_0_197), .ZN(n_0_0_193));
   INV_X1 i_0_0_352 (.A(n_0_0_194), .ZN(n_0_613));
   AOI221_X1 i_0_0_353 (.A(n_0_0_196), .B1(n_0_190), .B2(n_0_0_199), .C1(n_0_174), 
      .C2(n_0_0_198), .ZN(n_0_0_194));
   INV_X1 i_0_0_354 (.A(n_0_0_195), .ZN(n_0_614));
   AOI221_X1 i_0_0_355 (.A(n_0_0_196), .B1(n_0_191), .B2(n_0_0_199), .C1(n_0_175), 
      .C2(n_0_0_198), .ZN(n_0_0_195));
   AND2_X1 i_0_0_356 (.A1(n_0_629), .A2(n_0_0_197), .ZN(n_0_0_196));
   NOR2_X1 i_0_0_357 (.A1(n_0_0_199), .A2(n_0_0_198), .ZN(n_0_0_197));
   NOR2_X1 i_0_0_358 (.A1(n_0_0_333), .A2(multiplier[5]), .ZN(n_0_0_198));
   NOR2_X1 i_0_0_359 (.A1(multiplier[6]), .A2(n_0_0_332), .ZN(n_0_0_199));
   INV_X1 i_0_0_360 (.A(n_0_0_200), .ZN(product[5]));
   AOI222_X1 i_0_0_361 (.A1(n_0_128), .A2(n_0_0_218), .B1(n_0_144), .B2(
      n_0_0_219), .C1(n_0_630), .C2(n_0_0_217), .ZN(n_0_0_200));
   INV_X1 i_0_0_362 (.A(n_0_0_201), .ZN(n_0_615));
   AOI222_X1 i_0_0_363 (.A1(n_0_129), .A2(n_0_0_218), .B1(n_0_145), .B2(
      n_0_0_219), .C1(n_0_631), .C2(n_0_0_217), .ZN(n_0_0_201));
   INV_X1 i_0_0_364 (.A(n_0_0_202), .ZN(n_0_616));
   AOI222_X1 i_0_0_365 (.A1(n_0_130), .A2(n_0_0_218), .B1(n_0_146), .B2(
      n_0_0_219), .C1(n_0_632), .C2(n_0_0_217), .ZN(n_0_0_202));
   INV_X1 i_0_0_366 (.A(n_0_0_203), .ZN(n_0_617));
   AOI222_X1 i_0_0_367 (.A1(n_0_131), .A2(n_0_0_218), .B1(n_0_147), .B2(
      n_0_0_219), .C1(n_0_633), .C2(n_0_0_217), .ZN(n_0_0_203));
   INV_X1 i_0_0_368 (.A(n_0_0_204), .ZN(n_0_618));
   AOI222_X1 i_0_0_369 (.A1(n_0_132), .A2(n_0_0_218), .B1(n_0_148), .B2(
      n_0_0_219), .C1(n_0_634), .C2(n_0_0_217), .ZN(n_0_0_204));
   INV_X1 i_0_0_370 (.A(n_0_0_205), .ZN(n_0_619));
   AOI222_X1 i_0_0_371 (.A1(n_0_133), .A2(n_0_0_218), .B1(n_0_149), .B2(
      n_0_0_219), .C1(n_0_635), .C2(n_0_0_217), .ZN(n_0_0_205));
   INV_X1 i_0_0_372 (.A(n_0_0_206), .ZN(n_0_620));
   AOI222_X1 i_0_0_373 (.A1(n_0_134), .A2(n_0_0_218), .B1(n_0_150), .B2(
      n_0_0_219), .C1(n_0_636), .C2(n_0_0_217), .ZN(n_0_0_206));
   INV_X1 i_0_0_374 (.A(n_0_0_207), .ZN(n_0_621));
   AOI222_X1 i_0_0_375 (.A1(n_0_135), .A2(n_0_0_218), .B1(n_0_151), .B2(
      n_0_0_219), .C1(n_0_637), .C2(n_0_0_217), .ZN(n_0_0_207));
   INV_X1 i_0_0_376 (.A(n_0_0_208), .ZN(n_0_622));
   AOI222_X1 i_0_0_377 (.A1(n_0_136), .A2(n_0_0_218), .B1(n_0_152), .B2(
      n_0_0_219), .C1(n_0_638), .C2(n_0_0_217), .ZN(n_0_0_208));
   INV_X1 i_0_0_378 (.A(n_0_0_209), .ZN(n_0_623));
   AOI222_X1 i_0_0_379 (.A1(n_0_137), .A2(n_0_0_218), .B1(n_0_153), .B2(
      n_0_0_219), .C1(n_0_639), .C2(n_0_0_217), .ZN(n_0_0_209));
   INV_X1 i_0_0_380 (.A(n_0_0_210), .ZN(n_0_624));
   AOI222_X1 i_0_0_381 (.A1(n_0_154), .A2(n_0_0_219), .B1(n_0_138), .B2(
      n_0_0_218), .C1(n_0_640), .C2(n_0_0_217), .ZN(n_0_0_210));
   INV_X1 i_0_0_382 (.A(n_0_0_211), .ZN(n_0_625));
   AOI222_X1 i_0_0_383 (.A1(n_0_155), .A2(n_0_0_219), .B1(n_0_139), .B2(
      n_0_0_218), .C1(n_0_641), .C2(n_0_0_217), .ZN(n_0_0_211));
   INV_X1 i_0_0_384 (.A(n_0_0_212), .ZN(n_0_626));
   AOI222_X1 i_0_0_385 (.A1(n_0_156), .A2(n_0_0_219), .B1(n_0_140), .B2(
      n_0_0_218), .C1(n_0_642), .C2(n_0_0_217), .ZN(n_0_0_212));
   INV_X1 i_0_0_386 (.A(n_0_0_213), .ZN(n_0_627));
   AOI222_X1 i_0_0_387 (.A1(n_0_157), .A2(n_0_0_219), .B1(n_0_141), .B2(
      n_0_0_218), .C1(n_0_643), .C2(n_0_0_217), .ZN(n_0_0_213));
   INV_X1 i_0_0_388 (.A(n_0_0_214), .ZN(n_0_628));
   AOI221_X1 i_0_0_389 (.A(n_0_0_216), .B1(n_0_158), .B2(n_0_0_219), .C1(n_0_142), 
      .C2(n_0_0_218), .ZN(n_0_0_214));
   INV_X1 i_0_0_390 (.A(n_0_0_215), .ZN(n_0_629));
   AOI221_X1 i_0_0_391 (.A(n_0_0_216), .B1(n_0_159), .B2(n_0_0_219), .C1(n_0_143), 
      .C2(n_0_0_218), .ZN(n_0_0_215));
   AND2_X1 i_0_0_392 (.A1(n_0_644), .A2(n_0_0_217), .ZN(n_0_0_216));
   NOR2_X1 i_0_0_393 (.A1(n_0_0_219), .A2(n_0_0_218), .ZN(n_0_0_217));
   NOR2_X1 i_0_0_394 (.A1(n_0_0_332), .A2(multiplier[4]), .ZN(n_0_0_218));
   NOR2_X1 i_0_0_395 (.A1(multiplier[5]), .A2(n_0_0_331), .ZN(n_0_0_219));
   INV_X1 i_0_0_396 (.A(n_0_0_220), .ZN(product[4]));
   AOI222_X1 i_0_0_397 (.A1(n_0_96), .A2(n_0_0_238), .B1(n_0_112), .B2(n_0_0_239), 
      .C1(n_0_645), .C2(n_0_0_237), .ZN(n_0_0_220));
   INV_X1 i_0_0_398 (.A(n_0_0_221), .ZN(n_0_630));
   AOI222_X1 i_0_0_399 (.A1(n_0_97), .A2(n_0_0_238), .B1(n_0_113), .B2(n_0_0_239), 
      .C1(n_0_646), .C2(n_0_0_237), .ZN(n_0_0_221));
   INV_X1 i_0_0_400 (.A(n_0_0_222), .ZN(n_0_631));
   AOI222_X1 i_0_0_401 (.A1(n_0_98), .A2(n_0_0_238), .B1(n_0_114), .B2(n_0_0_239), 
      .C1(n_0_647), .C2(n_0_0_237), .ZN(n_0_0_222));
   INV_X1 i_0_0_402 (.A(n_0_0_223), .ZN(n_0_632));
   AOI222_X1 i_0_0_403 (.A1(n_0_99), .A2(n_0_0_238), .B1(n_0_115), .B2(n_0_0_239), 
      .C1(n_0_648), .C2(n_0_0_237), .ZN(n_0_0_223));
   INV_X1 i_0_0_404 (.A(n_0_0_224), .ZN(n_0_633));
   AOI222_X1 i_0_0_405 (.A1(n_0_100), .A2(n_0_0_238), .B1(n_0_116), .B2(
      n_0_0_239), .C1(n_0_649), .C2(n_0_0_237), .ZN(n_0_0_224));
   INV_X1 i_0_0_406 (.A(n_0_0_225), .ZN(n_0_634));
   AOI222_X1 i_0_0_407 (.A1(n_0_101), .A2(n_0_0_238), .B1(n_0_117), .B2(
      n_0_0_239), .C1(n_0_650), .C2(n_0_0_237), .ZN(n_0_0_225));
   INV_X1 i_0_0_408 (.A(n_0_0_226), .ZN(n_0_635));
   AOI222_X1 i_0_0_409 (.A1(n_0_102), .A2(n_0_0_238), .B1(n_0_118), .B2(
      n_0_0_239), .C1(n_0_651), .C2(n_0_0_237), .ZN(n_0_0_226));
   INV_X1 i_0_0_410 (.A(n_0_0_227), .ZN(n_0_636));
   AOI222_X1 i_0_0_411 (.A1(n_0_103), .A2(n_0_0_238), .B1(n_0_119), .B2(
      n_0_0_239), .C1(n_0_652), .C2(n_0_0_237), .ZN(n_0_0_227));
   INV_X1 i_0_0_412 (.A(n_0_0_228), .ZN(n_0_637));
   AOI222_X1 i_0_0_413 (.A1(n_0_104), .A2(n_0_0_238), .B1(n_0_120), .B2(
      n_0_0_239), .C1(n_0_653), .C2(n_0_0_237), .ZN(n_0_0_228));
   INV_X1 i_0_0_414 (.A(n_0_0_229), .ZN(n_0_638));
   AOI222_X1 i_0_0_415 (.A1(n_0_105), .A2(n_0_0_238), .B1(n_0_121), .B2(
      n_0_0_239), .C1(n_0_654), .C2(n_0_0_237), .ZN(n_0_0_229));
   INV_X1 i_0_0_416 (.A(n_0_0_230), .ZN(n_0_639));
   AOI222_X1 i_0_0_417 (.A1(n_0_106), .A2(n_0_0_238), .B1(n_0_122), .B2(
      n_0_0_239), .C1(n_0_655), .C2(n_0_0_237), .ZN(n_0_0_230));
   INV_X1 i_0_0_418 (.A(n_0_0_231), .ZN(n_0_640));
   AOI222_X1 i_0_0_419 (.A1(n_0_123), .A2(n_0_0_239), .B1(n_0_107), .B2(
      n_0_0_238), .C1(n_0_656), .C2(n_0_0_237), .ZN(n_0_0_231));
   INV_X1 i_0_0_420 (.A(n_0_0_232), .ZN(n_0_641));
   AOI222_X1 i_0_0_421 (.A1(n_0_124), .A2(n_0_0_239), .B1(n_0_108), .B2(
      n_0_0_238), .C1(n_0_657), .C2(n_0_0_237), .ZN(n_0_0_232));
   INV_X1 i_0_0_422 (.A(n_0_0_233), .ZN(n_0_642));
   AOI222_X1 i_0_0_423 (.A1(n_0_125), .A2(n_0_0_239), .B1(n_0_109), .B2(
      n_0_0_238), .C1(n_0_658), .C2(n_0_0_237), .ZN(n_0_0_233));
   INV_X1 i_0_0_424 (.A(n_0_0_234), .ZN(n_0_643));
   AOI221_X1 i_0_0_425 (.A(n_0_0_236), .B1(n_0_126), .B2(n_0_0_239), .C1(n_0_110), 
      .C2(n_0_0_238), .ZN(n_0_0_234));
   INV_X1 i_0_0_426 (.A(n_0_0_235), .ZN(n_0_644));
   AOI221_X1 i_0_0_427 (.A(n_0_0_236), .B1(n_0_127), .B2(n_0_0_239), .C1(n_0_111), 
      .C2(n_0_0_238), .ZN(n_0_0_235));
   AND2_X1 i_0_0_428 (.A1(n_0_659), .A2(n_0_0_237), .ZN(n_0_0_236));
   NOR2_X1 i_0_0_429 (.A1(n_0_0_239), .A2(n_0_0_238), .ZN(n_0_0_237));
   NOR2_X1 i_0_0_430 (.A1(n_0_0_331), .A2(multiplier[3]), .ZN(n_0_0_238));
   NOR2_X1 i_0_0_431 (.A1(multiplier[4]), .A2(n_0_0_330), .ZN(n_0_0_239));
   INV_X1 i_0_0_432 (.A(n_0_0_240), .ZN(product[3]));
   AOI222_X1 i_0_0_433 (.A1(n_0_80), .A2(n_0_0_258), .B1(n_0_64), .B2(n_0_0_259), 
      .C1(n_0_660), .C2(n_0_0_257), .ZN(n_0_0_240));
   INV_X1 i_0_0_434 (.A(n_0_0_241), .ZN(n_0_645));
   AOI222_X1 i_0_0_435 (.A1(n_0_81), .A2(n_0_0_258), .B1(n_0_65), .B2(n_0_0_259), 
      .C1(n_0_661), .C2(n_0_0_257), .ZN(n_0_0_241));
   INV_X1 i_0_0_436 (.A(n_0_0_242), .ZN(n_0_646));
   AOI222_X1 i_0_0_437 (.A1(n_0_82), .A2(n_0_0_258), .B1(n_0_66), .B2(n_0_0_259), 
      .C1(n_0_662), .C2(n_0_0_257), .ZN(n_0_0_242));
   INV_X1 i_0_0_438 (.A(n_0_0_243), .ZN(n_0_647));
   AOI222_X1 i_0_0_439 (.A1(n_0_83), .A2(n_0_0_258), .B1(n_0_67), .B2(n_0_0_259), 
      .C1(n_0_663), .C2(n_0_0_257), .ZN(n_0_0_243));
   INV_X1 i_0_0_440 (.A(n_0_0_244), .ZN(n_0_648));
   AOI222_X1 i_0_0_441 (.A1(n_0_84), .A2(n_0_0_258), .B1(n_0_68), .B2(n_0_0_259), 
      .C1(n_0_664), .C2(n_0_0_257), .ZN(n_0_0_244));
   INV_X1 i_0_0_442 (.A(n_0_0_245), .ZN(n_0_649));
   AOI222_X1 i_0_0_443 (.A1(n_0_85), .A2(n_0_0_258), .B1(n_0_69), .B2(n_0_0_259), 
      .C1(n_0_665), .C2(n_0_0_257), .ZN(n_0_0_245));
   INV_X1 i_0_0_444 (.A(n_0_0_246), .ZN(n_0_650));
   AOI222_X1 i_0_0_445 (.A1(n_0_86), .A2(n_0_0_258), .B1(n_0_70), .B2(n_0_0_259), 
      .C1(n_0_666), .C2(n_0_0_257), .ZN(n_0_0_246));
   INV_X1 i_0_0_446 (.A(n_0_0_247), .ZN(n_0_651));
   AOI222_X1 i_0_0_447 (.A1(n_0_87), .A2(n_0_0_258), .B1(n_0_71), .B2(n_0_0_259), 
      .C1(n_0_667), .C2(n_0_0_257), .ZN(n_0_0_247));
   INV_X1 i_0_0_448 (.A(n_0_0_248), .ZN(n_0_652));
   AOI222_X1 i_0_0_449 (.A1(n_0_88), .A2(n_0_0_258), .B1(n_0_72), .B2(n_0_0_259), 
      .C1(n_0_668), .C2(n_0_0_257), .ZN(n_0_0_248));
   INV_X1 i_0_0_450 (.A(n_0_0_249), .ZN(n_0_653));
   AOI222_X1 i_0_0_451 (.A1(n_0_89), .A2(n_0_0_258), .B1(n_0_73), .B2(n_0_0_259), 
      .C1(n_0_669), .C2(n_0_0_257), .ZN(n_0_0_249));
   INV_X1 i_0_0_452 (.A(n_0_0_250), .ZN(n_0_654));
   AOI222_X1 i_0_0_453 (.A1(n_0_90), .A2(n_0_0_258), .B1(n_0_74), .B2(n_0_0_259), 
      .C1(n_0_670), .C2(n_0_0_257), .ZN(n_0_0_250));
   INV_X1 i_0_0_454 (.A(n_0_0_251), .ZN(n_0_655));
   AOI222_X1 i_0_0_455 (.A1(n_0_91), .A2(n_0_0_258), .B1(n_0_75), .B2(n_0_0_259), 
      .C1(n_0_671), .C2(n_0_0_257), .ZN(n_0_0_251));
   INV_X1 i_0_0_456 (.A(n_0_0_252), .ZN(n_0_656));
   AOI222_X1 i_0_0_457 (.A1(n_0_76), .A2(n_0_0_259), .B1(n_0_92), .B2(n_0_0_258), 
      .C1(n_0_672), .C2(n_0_0_257), .ZN(n_0_0_252));
   INV_X1 i_0_0_458 (.A(n_0_0_253), .ZN(n_0_657));
   AOI222_X1 i_0_0_459 (.A1(n_0_77), .A2(n_0_0_259), .B1(n_0_93), .B2(n_0_0_258), 
      .C1(n_0_673), .C2(n_0_0_257), .ZN(n_0_0_253));
   INV_X1 i_0_0_460 (.A(n_0_0_254), .ZN(n_0_658));
   AOI221_X1 i_0_0_461 (.A(n_0_0_256), .B1(n_0_78), .B2(n_0_0_259), .C1(n_0_94), 
      .C2(n_0_0_258), .ZN(n_0_0_254));
   INV_X1 i_0_0_462 (.A(n_0_0_255), .ZN(n_0_659));
   AOI221_X1 i_0_0_463 (.A(n_0_0_256), .B1(n_0_79), .B2(n_0_0_259), .C1(n_0_95), 
      .C2(n_0_0_258), .ZN(n_0_0_255));
   AND2_X1 i_0_0_464 (.A1(n_0_674), .A2(n_0_0_257), .ZN(n_0_0_256));
   NOR2_X1 i_0_0_465 (.A1(n_0_0_259), .A2(n_0_0_258), .ZN(n_0_0_257));
   NOR2_X1 i_0_0_466 (.A1(multiplier[3]), .A2(n_0_0_329), .ZN(n_0_0_258));
   NOR2_X1 i_0_0_467 (.A1(n_0_0_330), .A2(multiplier[2]), .ZN(n_0_0_259));
   INV_X1 i_0_0_468 (.A(n_0_0_260), .ZN(product[2]));
   AOI222_X1 i_0_0_469 (.A1(n_0_32), .A2(n_0_0_278), .B1(n_0_48), .B2(n_0_0_279), 
      .C1(n_0_675), .C2(n_0_0_277), .ZN(n_0_0_260));
   INV_X1 i_0_0_470 (.A(n_0_0_261), .ZN(n_0_660));
   AOI222_X1 i_0_0_471 (.A1(n_0_33), .A2(n_0_0_278), .B1(n_0_49), .B2(n_0_0_279), 
      .C1(n_0_676), .C2(n_0_0_277), .ZN(n_0_0_261));
   INV_X1 i_0_0_472 (.A(n_0_0_262), .ZN(n_0_661));
   AOI222_X1 i_0_0_473 (.A1(n_0_34), .A2(n_0_0_278), .B1(n_0_50), .B2(n_0_0_279), 
      .C1(n_0_677), .C2(n_0_0_277), .ZN(n_0_0_262));
   INV_X1 i_0_0_474 (.A(n_0_0_263), .ZN(n_0_662));
   AOI222_X1 i_0_0_475 (.A1(n_0_35), .A2(n_0_0_278), .B1(n_0_51), .B2(n_0_0_279), 
      .C1(n_0_678), .C2(n_0_0_277), .ZN(n_0_0_263));
   INV_X1 i_0_0_476 (.A(n_0_0_264), .ZN(n_0_663));
   AOI222_X1 i_0_0_477 (.A1(n_0_36), .A2(n_0_0_278), .B1(n_0_52), .B2(n_0_0_279), 
      .C1(n_0_679), .C2(n_0_0_277), .ZN(n_0_0_264));
   INV_X1 i_0_0_478 (.A(n_0_0_265), .ZN(n_0_664));
   AOI222_X1 i_0_0_479 (.A1(n_0_37), .A2(n_0_0_278), .B1(n_0_53), .B2(n_0_0_279), 
      .C1(n_0_680), .C2(n_0_0_277), .ZN(n_0_0_265));
   INV_X1 i_0_0_480 (.A(n_0_0_266), .ZN(n_0_665));
   AOI222_X1 i_0_0_481 (.A1(n_0_38), .A2(n_0_0_278), .B1(n_0_54), .B2(n_0_0_279), 
      .C1(n_0_681), .C2(n_0_0_277), .ZN(n_0_0_266));
   INV_X1 i_0_0_482 (.A(n_0_0_267), .ZN(n_0_666));
   AOI222_X1 i_0_0_483 (.A1(n_0_39), .A2(n_0_0_278), .B1(n_0_55), .B2(n_0_0_279), 
      .C1(n_0_682), .C2(n_0_0_277), .ZN(n_0_0_267));
   INV_X1 i_0_0_484 (.A(n_0_0_268), .ZN(n_0_667));
   AOI222_X1 i_0_0_485 (.A1(n_0_40), .A2(n_0_0_278), .B1(n_0_56), .B2(n_0_0_279), 
      .C1(n_0_683), .C2(n_0_0_277), .ZN(n_0_0_268));
   INV_X1 i_0_0_486 (.A(n_0_0_269), .ZN(n_0_668));
   AOI222_X1 i_0_0_487 (.A1(n_0_41), .A2(n_0_0_278), .B1(n_0_57), .B2(n_0_0_279), 
      .C1(n_0_684), .C2(n_0_0_277), .ZN(n_0_0_269));
   INV_X1 i_0_0_488 (.A(n_0_0_270), .ZN(n_0_669));
   AOI222_X1 i_0_0_489 (.A1(n_0_42), .A2(n_0_0_278), .B1(n_0_58), .B2(n_0_0_279), 
      .C1(n_0_685), .C2(n_0_0_277), .ZN(n_0_0_270));
   INV_X1 i_0_0_490 (.A(n_0_0_271), .ZN(n_0_670));
   AOI222_X1 i_0_0_491 (.A1(n_0_59), .A2(n_0_0_279), .B1(n_0_43), .B2(n_0_0_278), 
      .C1(n_0_686), .C2(n_0_0_277), .ZN(n_0_0_271));
   INV_X1 i_0_0_492 (.A(n_0_0_272), .ZN(n_0_671));
   AOI222_X1 i_0_0_493 (.A1(n_0_44), .A2(n_0_0_278), .B1(n_0_60), .B2(n_0_0_279), 
      .C1(n_0_687), .C2(n_0_0_277), .ZN(n_0_0_272));
   INV_X1 i_0_0_494 (.A(n_0_0_273), .ZN(n_0_672));
   AOI222_X1 i_0_0_495 (.A1(n_0_45), .A2(n_0_0_278), .B1(n_0_61), .B2(n_0_0_279), 
      .C1(n_0_688), .C2(n_0_0_277), .ZN(n_0_0_273));
   INV_X1 i_0_0_496 (.A(n_0_0_274), .ZN(n_0_673));
   AOI221_X1 i_0_0_497 (.A(n_0_0_276), .B1(n_0_62), .B2(n_0_0_279), .C1(n_0_46), 
      .C2(n_0_0_278), .ZN(n_0_0_274));
   INV_X1 i_0_0_498 (.A(n_0_0_275), .ZN(n_0_674));
   AOI221_X1 i_0_0_499 (.A(n_0_0_276), .B1(n_0_63), .B2(n_0_0_279), .C1(n_0_47), 
      .C2(n_0_0_278), .ZN(n_0_0_275));
   AND2_X1 i_0_0_500 (.A1(n_0_689), .A2(n_0_0_277), .ZN(n_0_0_276));
   NOR2_X1 i_0_0_501 (.A1(n_0_0_279), .A2(n_0_0_278), .ZN(n_0_0_277));
   NOR2_X1 i_0_0_502 (.A1(n_0_0_329), .A2(multiplier[1]), .ZN(n_0_0_278));
   NOR2_X1 i_0_0_503 (.A1(multiplier[2]), .A2(n_0_0_328), .ZN(n_0_0_279));
   INV_X1 i_0_0_504 (.A(n_0_0_280), .ZN(product[1]));
   AOI222_X1 i_0_0_505 (.A1(n_0_16), .A2(n_0_0_296), .B1(n_0_0), .B2(n_0_0_297), 
      .C1(n_0_705), .C2(n_0_0_299), .ZN(n_0_0_280));
   INV_X1 i_0_0_506 (.A(n_0_0_281), .ZN(n_0_675));
   AOI222_X1 i_0_0_507 (.A1(n_0_17), .A2(n_0_0_296), .B1(n_0_1), .B2(n_0_0_297), 
      .C1(n_0_706), .C2(n_0_0_299), .ZN(n_0_0_281));
   INV_X1 i_0_0_508 (.A(n_0_0_282), .ZN(n_0_676));
   AOI222_X1 i_0_0_509 (.A1(n_0_18), .A2(n_0_0_296), .B1(n_0_2), .B2(n_0_0_297), 
      .C1(n_0_707), .C2(n_0_0_299), .ZN(n_0_0_282));
   INV_X1 i_0_0_510 (.A(n_0_0_283), .ZN(n_0_677));
   AOI222_X1 i_0_0_511 (.A1(n_0_19), .A2(n_0_0_296), .B1(n_0_3), .B2(n_0_0_297), 
      .C1(n_0_708), .C2(n_0_0_299), .ZN(n_0_0_283));
   INV_X1 i_0_0_512 (.A(n_0_0_284), .ZN(n_0_678));
   AOI222_X1 i_0_0_513 (.A1(n_0_20), .A2(n_0_0_296), .B1(n_0_4), .B2(n_0_0_297), 
      .C1(n_0_709), .C2(n_0_0_299), .ZN(n_0_0_284));
   INV_X1 i_0_0_514 (.A(n_0_0_285), .ZN(n_0_679));
   AOI222_X1 i_0_0_515 (.A1(n_0_21), .A2(n_0_0_296), .B1(n_0_5), .B2(n_0_0_297), 
      .C1(n_0_710), .C2(n_0_0_299), .ZN(n_0_0_285));
   INV_X1 i_0_0_516 (.A(n_0_0_286), .ZN(n_0_680));
   AOI222_X1 i_0_0_517 (.A1(n_0_22), .A2(n_0_0_296), .B1(n_0_6), .B2(n_0_0_297), 
      .C1(n_0_711), .C2(n_0_0_299), .ZN(n_0_0_286));
   INV_X1 i_0_0_518 (.A(n_0_0_287), .ZN(n_0_681));
   AOI222_X1 i_0_0_519 (.A1(n_0_23), .A2(n_0_0_296), .B1(n_0_7), .B2(n_0_0_297), 
      .C1(n_0_712), .C2(n_0_0_299), .ZN(n_0_0_287));
   INV_X1 i_0_0_520 (.A(n_0_0_288), .ZN(n_0_682));
   AOI222_X1 i_0_0_521 (.A1(n_0_24), .A2(n_0_0_296), .B1(n_0_8), .B2(n_0_0_297), 
      .C1(n_0_713), .C2(n_0_0_299), .ZN(n_0_0_288));
   INV_X1 i_0_0_522 (.A(n_0_0_289), .ZN(n_0_683));
   AOI222_X1 i_0_0_523 (.A1(n_0_25), .A2(n_0_0_296), .B1(n_0_9), .B2(n_0_0_297), 
      .C1(n_0_714), .C2(n_0_0_299), .ZN(n_0_0_289));
   INV_X1 i_0_0_524 (.A(n_0_0_290), .ZN(n_0_684));
   AOI222_X1 i_0_0_525 (.A1(n_0_26), .A2(n_0_0_296), .B1(n_0_10), .B2(n_0_0_297), 
      .C1(n_0_715), .C2(n_0_0_299), .ZN(n_0_0_290));
   INV_X1 i_0_0_526 (.A(n_0_0_291), .ZN(n_0_685));
   AOI222_X1 i_0_0_527 (.A1(n_0_27), .A2(n_0_0_296), .B1(n_0_11), .B2(n_0_0_297), 
      .C1(n_0_716), .C2(n_0_0_299), .ZN(n_0_0_291));
   INV_X1 i_0_0_528 (.A(n_0_0_292), .ZN(n_0_686));
   AOI222_X1 i_0_0_529 (.A1(n_0_28), .A2(n_0_0_296), .B1(n_0_12), .B2(n_0_0_297), 
      .C1(n_0_717), .C2(n_0_0_299), .ZN(n_0_0_292));
   INV_X1 i_0_0_530 (.A(n_0_0_293), .ZN(n_0_687));
   AOI222_X1 i_0_0_531 (.A1(n_0_29), .A2(n_0_0_296), .B1(n_0_13), .B2(n_0_0_297), 
      .C1(n_0_718), .C2(n_0_0_299), .ZN(n_0_0_293));
   INV_X1 i_0_0_532 (.A(n_0_0_294), .ZN(n_0_688));
   AOI221_X1 i_0_0_533 (.A(n_0_0_298), .B1(n_0_30), .B2(n_0_0_296), .C1(n_0_14), 
      .C2(n_0_0_297), .ZN(n_0_0_294));
   INV_X1 i_0_0_534 (.A(n_0_0_295), .ZN(n_0_689));
   AOI221_X1 i_0_0_535 (.A(n_0_0_298), .B1(n_0_31), .B2(n_0_0_296), .C1(n_0_15), 
      .C2(n_0_0_297), .ZN(n_0_0_295));
   NOR2_X1 i_0_0_536 (.A1(multiplier[1]), .A2(n_0_0_327), .ZN(n_0_0_296));
   NOR2_X1 i_0_0_537 (.A1(n_0_0_328), .A2(multiplier[0]), .ZN(n_0_0_297));
   AND2_X1 i_0_0_538 (.A1(multiplier[1]), .A2(n_0_704), .ZN(n_0_0_298));
   NOR2_X1 i_0_0_539 (.A1(n_0_0_328), .A2(n_0_0_327), .ZN(n_0_0_299));
   AND2_X1 i_0_0_540 (.A1(multiplicand[0]), .A2(multiplier[0]), .ZN(product[0]));
   AND2_X1 i_0_0_541 (.A1(multiplier[0]), .A2(n_0_705), .ZN(n_0_690));
   AND2_X1 i_0_0_542 (.A1(multiplier[0]), .A2(n_0_706), .ZN(n_0_691));
   AND2_X1 i_0_0_543 (.A1(multiplier[0]), .A2(n_0_707), .ZN(n_0_692));
   AND2_X1 i_0_0_544 (.A1(multiplier[0]), .A2(n_0_708), .ZN(n_0_693));
   AND2_X1 i_0_0_545 (.A1(multiplier[0]), .A2(n_0_709), .ZN(n_0_694));
   AND2_X1 i_0_0_546 (.A1(multiplier[0]), .A2(n_0_710), .ZN(n_0_695));
   AND2_X1 i_0_0_547 (.A1(multiplier[0]), .A2(n_0_711), .ZN(n_0_696));
   AND2_X1 i_0_0_548 (.A1(multiplier[0]), .A2(n_0_712), .ZN(n_0_697));
   AND2_X1 i_0_0_549 (.A1(multiplier[0]), .A2(n_0_713), .ZN(n_0_698));
   AND2_X1 i_0_0_550 (.A1(multiplier[0]), .A2(n_0_714), .ZN(n_0_699));
   AND2_X1 i_0_0_551 (.A1(multiplier[0]), .A2(n_0_715), .ZN(n_0_700));
   AND2_X1 i_0_0_552 (.A1(multiplier[0]), .A2(n_0_716), .ZN(n_0_701));
   AND2_X1 i_0_0_553 (.A1(multiplier[0]), .A2(n_0_717), .ZN(n_0_702));
   AND2_X1 i_0_0_554 (.A1(multiplier[0]), .A2(n_0_718), .ZN(n_0_703));
   AND2_X1 i_0_0_555 (.A1(multiplier[0]), .A2(n_0_719), .ZN(n_0_704));
   AOI21_X1 i_0_0_556 (.A(n_0_0_326), .B1(multiplicand[1]), .B2(multiplicand[0]), 
      .ZN(n_0_705));
   AOI21_X1 i_0_0_557 (.A(n_0_0_324), .B1(multiplicand[2]), .B2(n_0_0_325), 
      .ZN(n_0_706));
   AOI21_X1 i_0_0_558 (.A(n_0_0_322), .B1(multiplicand[3]), .B2(n_0_0_323), 
      .ZN(n_0_707));
   AOI21_X1 i_0_0_559 (.A(n_0_0_320), .B1(multiplicand[4]), .B2(n_0_0_321), 
      .ZN(n_0_708));
   AOI21_X1 i_0_0_560 (.A(n_0_0_318), .B1(multiplicand[5]), .B2(n_0_0_319), 
      .ZN(n_0_709));
   AOI21_X1 i_0_0_561 (.A(n_0_0_316), .B1(multiplicand[6]), .B2(n_0_0_317), 
      .ZN(n_0_710));
   AOI21_X1 i_0_0_562 (.A(n_0_0_314), .B1(multiplicand[7]), .B2(n_0_0_315), 
      .ZN(n_0_711));
   AOI21_X1 i_0_0_563 (.A(n_0_0_312), .B1(multiplicand[8]), .B2(n_0_0_313), 
      .ZN(n_0_712));
   AOI21_X1 i_0_0_564 (.A(n_0_0_310), .B1(multiplicand[9]), .B2(n_0_0_311), 
      .ZN(n_0_713));
   AOI21_X1 i_0_0_565 (.A(n_0_0_308), .B1(multiplicand[10]), .B2(n_0_0_309), 
      .ZN(n_0_714));
   AOI21_X1 i_0_0_566 (.A(n_0_0_306), .B1(multiplicand[11]), .B2(n_0_0_307), 
      .ZN(n_0_715));
   AOI21_X1 i_0_0_567 (.A(n_0_0_304), .B1(multiplicand[12]), .B2(n_0_0_305), 
      .ZN(n_0_716));
   AOI21_X1 i_0_0_568 (.A(n_0_0_302), .B1(multiplicand[13]), .B2(n_0_0_303), 
      .ZN(n_0_717));
   AOI21_X1 i_0_0_569 (.A(n_0_0_300), .B1(multiplicand[14]), .B2(n_0_0_301), 
      .ZN(n_0_718));
   XNOR2_X1 i_0_0_570 (.A(multiplicand[15]), .B(n_0_0_300), .ZN(n_0_719));
   NOR2_X1 i_0_0_571 (.A1(multiplicand[14]), .A2(n_0_0_301), .ZN(n_0_0_300));
   INV_X1 i_0_0_572 (.A(n_0_0_302), .ZN(n_0_0_301));
   NOR2_X1 i_0_0_573 (.A1(multiplicand[13]), .A2(n_0_0_303), .ZN(n_0_0_302));
   INV_X1 i_0_0_574 (.A(n_0_0_304), .ZN(n_0_0_303));
   NOR2_X1 i_0_0_575 (.A1(multiplicand[12]), .A2(n_0_0_305), .ZN(n_0_0_304));
   INV_X1 i_0_0_576 (.A(n_0_0_306), .ZN(n_0_0_305));
   NOR2_X1 i_0_0_577 (.A1(multiplicand[11]), .A2(n_0_0_307), .ZN(n_0_0_306));
   INV_X1 i_0_0_578 (.A(n_0_0_308), .ZN(n_0_0_307));
   NOR2_X1 i_0_0_579 (.A1(multiplicand[10]), .A2(n_0_0_309), .ZN(n_0_0_308));
   INV_X1 i_0_0_580 (.A(n_0_0_310), .ZN(n_0_0_309));
   NOR2_X1 i_0_0_581 (.A1(multiplicand[9]), .A2(n_0_0_311), .ZN(n_0_0_310));
   INV_X1 i_0_0_582 (.A(n_0_0_312), .ZN(n_0_0_311));
   NOR2_X1 i_0_0_583 (.A1(multiplicand[8]), .A2(n_0_0_313), .ZN(n_0_0_312));
   INV_X1 i_0_0_584 (.A(n_0_0_314), .ZN(n_0_0_313));
   NOR2_X1 i_0_0_585 (.A1(multiplicand[7]), .A2(n_0_0_315), .ZN(n_0_0_314));
   INV_X1 i_0_0_586 (.A(n_0_0_316), .ZN(n_0_0_315));
   NOR2_X1 i_0_0_587 (.A1(multiplicand[6]), .A2(n_0_0_317), .ZN(n_0_0_316));
   INV_X1 i_0_0_588 (.A(n_0_0_318), .ZN(n_0_0_317));
   NOR2_X1 i_0_0_589 (.A1(multiplicand[5]), .A2(n_0_0_319), .ZN(n_0_0_318));
   INV_X1 i_0_0_590 (.A(n_0_0_320), .ZN(n_0_0_319));
   NOR2_X1 i_0_0_591 (.A1(multiplicand[4]), .A2(n_0_0_321), .ZN(n_0_0_320));
   INV_X1 i_0_0_592 (.A(n_0_0_322), .ZN(n_0_0_321));
   NOR2_X1 i_0_0_593 (.A1(multiplicand[3]), .A2(n_0_0_323), .ZN(n_0_0_322));
   INV_X1 i_0_0_594 (.A(n_0_0_324), .ZN(n_0_0_323));
   NOR2_X1 i_0_0_595 (.A1(multiplicand[2]), .A2(n_0_0_325), .ZN(n_0_0_324));
   INV_X1 i_0_0_596 (.A(n_0_0_326), .ZN(n_0_0_325));
   NOR2_X1 i_0_0_597 (.A1(multiplicand[1]), .A2(multiplicand[0]), .ZN(n_0_0_326));
   INV_X1 i_0_0_598 (.A(multiplier[0]), .ZN(n_0_0_327));
   INV_X1 i_0_0_599 (.A(multiplier[1]), .ZN(n_0_0_328));
   INV_X1 i_0_0_600 (.A(multiplier[2]), .ZN(n_0_0_329));
   INV_X1 i_0_0_601 (.A(multiplier[3]), .ZN(n_0_0_330));
   INV_X1 i_0_0_602 (.A(multiplier[4]), .ZN(n_0_0_331));
   INV_X1 i_0_0_603 (.A(multiplier[5]), .ZN(n_0_0_332));
   INV_X1 i_0_0_604 (.A(multiplier[6]), .ZN(n_0_0_333));
   INV_X1 i_0_0_605 (.A(multiplier[7]), .ZN(n_0_0_334));
   INV_X1 i_0_0_606 (.A(multiplier[8]), .ZN(n_0_0_335));
   INV_X1 i_0_0_607 (.A(multiplier[9]), .ZN(n_0_0_336));
   INV_X1 i_0_0_608 (.A(multiplier[10]), .ZN(n_0_0_337));
   INV_X1 i_0_0_609 (.A(multiplier[11]), .ZN(n_0_0_338));
   INV_X1 i_0_0_610 (.A(multiplier[12]), .ZN(n_0_0_339));
   INV_X1 i_0_0_611 (.A(multiplier[13]), .ZN(n_0_0_340));
   INV_X1 i_0_0_612 (.A(multiplier[14]), .ZN(n_0_0_341));
endmodule
