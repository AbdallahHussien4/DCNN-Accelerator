/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Wed May 26 02:27:45 2021
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 2140351355 */

module RAM(enable, clk, address, write, \output_data[0][0] , \output_data[0][1] , 
      \output_data[0][2] , \output_data[0][3] , \output_data[0][4] , 
      \output_data[1][0] , \output_data[1][1] , \output_data[1][2] , 
      \output_data[1][3] , \output_data[1][4] , \output_data[2][0] , 
      \output_data[2][1] , \output_data[2][2] , \output_data[2][3] , 
      \output_data[2][4] , \output_data[3][0] , \output_data[3][1] , 
      \output_data[3][2] , \output_data[3][3] , \output_data[3][4] , 
      \output_data[4][0] , \output_data[4][1] , \output_data[4][2] , 
      \output_data[4][3] , \output_data[4][4] , offset, input_data, finish);
   input enable;
   input clk;
   input [15:0]address;
   input write;
   output [15:0]\output_data[0][0] ;
   output [15:0]\output_data[0][1] ;
   output [15:0]\output_data[0][2] ;
   output [15:0]\output_data[0][3] ;
   output [15:0]\output_data[0][4] ;
   output [15:0]\output_data[1][0] ;
   output [15:0]\output_data[1][1] ;
   output [15:0]\output_data[1][2] ;
   output [15:0]\output_data[1][3] ;
   output [15:0]\output_data[1][4] ;
   output [15:0]\output_data[2][0] ;
   output [15:0]\output_data[2][1] ;
   output [15:0]\output_data[2][2] ;
   output [15:0]\output_data[2][3] ;
   output [15:0]\output_data[2][4] ;
   output [15:0]\output_data[3][0] ;
   output [15:0]\output_data[3][1] ;
   output [15:0]\output_data[3][2] ;
   output [15:0]\output_data[3][3] ;
   output [15:0]\output_data[3][4] ;
   output [15:0]\output_data[4][0] ;
   output [15:0]\output_data[4][1] ;
   output [15:0]\output_data[4][2] ;
   output [15:0]\output_data[4][3] ;
   output [15:0]\output_data[4][4] ;
   input [15:0]offset;
   input [15:0]input_data;
   output finish;

   wire n_27_0;

   assign \output_data[0][0] [15] = 1'b0;
   assign \output_data[0][0] [14] = 1'b0;
   assign \output_data[0][0] [13] = 1'b0;
   assign \output_data[0][0] [12] = 1'b0;
   assign \output_data[0][0] [11] = 1'b0;
   assign \output_data[0][0] [10] = 1'b0;
   assign \output_data[0][0] [9] = 1'b0;
   assign \output_data[0][0] [8] = 1'b0;
   assign \output_data[0][0] [7] = 1'b0;
   assign \output_data[0][0] [6] = 1'b0;
   assign \output_data[0][0] [5] = 1'b0;
   assign \output_data[0][0] [4] = 1'b0;
   assign \output_data[0][0] [3] = 1'b0;
   assign \output_data[0][0] [2] = 1'b0;
   assign \output_data[0][0] [1] = 1'b0;
   assign \output_data[0][0] [0] = 1'b0;
   assign \output_data[0][1] [15] = 1'b0;
   assign \output_data[0][1] [14] = 1'b0;
   assign \output_data[0][1] [13] = 1'b0;
   assign \output_data[0][1] [12] = 1'b0;
   assign \output_data[0][1] [11] = 1'b0;
   assign \output_data[0][1] [10] = 1'b0;
   assign \output_data[0][1] [9] = 1'b0;
   assign \output_data[0][1] [8] = 1'b0;
   assign \output_data[0][1] [7] = 1'b0;
   assign \output_data[0][1] [6] = 1'b0;
   assign \output_data[0][1] [5] = 1'b0;
   assign \output_data[0][1] [4] = 1'b0;
   assign \output_data[0][1] [3] = 1'b0;
   assign \output_data[0][1] [2] = 1'b0;
   assign \output_data[0][1] [1] = 1'b0;
   assign \output_data[0][1] [0] = 1'b0;
   assign \output_data[0][2] [15] = 1'b0;
   assign \output_data[0][2] [14] = 1'b0;
   assign \output_data[0][2] [13] = 1'b0;
   assign \output_data[0][2] [12] = 1'b0;
   assign \output_data[0][2] [11] = 1'b0;
   assign \output_data[0][2] [10] = 1'b0;
   assign \output_data[0][2] [9] = 1'b0;
   assign \output_data[0][2] [8] = 1'b0;
   assign \output_data[0][2] [7] = 1'b0;
   assign \output_data[0][2] [6] = 1'b0;
   assign \output_data[0][2] [5] = 1'b0;
   assign \output_data[0][2] [4] = 1'b0;
   assign \output_data[0][2] [3] = 1'b0;
   assign \output_data[0][2] [2] = 1'b0;
   assign \output_data[0][2] [1] = 1'b0;
   assign \output_data[0][2] [0] = 1'b0;
   assign \output_data[0][3] [15] = 1'b0;
   assign \output_data[0][3] [14] = 1'b0;
   assign \output_data[0][3] [13] = 1'b0;
   assign \output_data[0][3] [12] = 1'b0;
   assign \output_data[0][3] [11] = 1'b0;
   assign \output_data[0][3] [10] = 1'b0;
   assign \output_data[0][3] [9] = 1'b0;
   assign \output_data[0][3] [8] = 1'b0;
   assign \output_data[0][3] [7] = 1'b0;
   assign \output_data[0][3] [6] = 1'b0;
   assign \output_data[0][3] [5] = 1'b0;
   assign \output_data[0][3] [4] = 1'b0;
   assign \output_data[0][3] [3] = 1'b0;
   assign \output_data[0][3] [2] = 1'b0;
   assign \output_data[0][3] [1] = 1'b0;
   assign \output_data[0][3] [0] = 1'b0;
   assign \output_data[0][4] [15] = 1'b0;
   assign \output_data[0][4] [14] = 1'b0;
   assign \output_data[0][4] [13] = 1'b0;
   assign \output_data[0][4] [12] = 1'b0;
   assign \output_data[0][4] [11] = 1'b0;
   assign \output_data[0][4] [10] = 1'b0;
   assign \output_data[0][4] [9] = 1'b0;
   assign \output_data[0][4] [8] = 1'b0;
   assign \output_data[0][4] [7] = 1'b0;
   assign \output_data[0][4] [6] = 1'b0;
   assign \output_data[0][4] [5] = 1'b0;
   assign \output_data[0][4] [4] = 1'b0;
   assign \output_data[0][4] [3] = 1'b0;
   assign \output_data[0][4] [2] = 1'b0;
   assign \output_data[0][4] [1] = 1'b0;
   assign \output_data[0][4] [0] = 1'b0;
   assign \output_data[1][0] [15] = 1'b0;
   assign \output_data[1][0] [14] = 1'b0;
   assign \output_data[1][0] [13] = 1'b0;
   assign \output_data[1][0] [12] = 1'b0;
   assign \output_data[1][0] [11] = 1'b0;
   assign \output_data[1][0] [10] = 1'b0;
   assign \output_data[1][0] [9] = 1'b0;
   assign \output_data[1][0] [8] = 1'b0;
   assign \output_data[1][0] [7] = 1'b0;
   assign \output_data[1][0] [6] = 1'b0;
   assign \output_data[1][0] [5] = 1'b0;
   assign \output_data[1][0] [4] = 1'b0;
   assign \output_data[1][0] [3] = 1'b0;
   assign \output_data[1][0] [2] = 1'b0;
   assign \output_data[1][0] [1] = 1'b0;
   assign \output_data[1][0] [0] = 1'b0;
   assign \output_data[1][1] [15] = 1'b0;
   assign \output_data[1][1] [14] = 1'b0;
   assign \output_data[1][1] [13] = 1'b0;
   assign \output_data[1][1] [12] = 1'b0;
   assign \output_data[1][1] [11] = 1'b0;
   assign \output_data[1][1] [10] = 1'b0;
   assign \output_data[1][1] [9] = 1'b0;
   assign \output_data[1][1] [8] = 1'b0;
   assign \output_data[1][1] [7] = 1'b0;
   assign \output_data[1][1] [6] = 1'b0;
   assign \output_data[1][1] [5] = 1'b0;
   assign \output_data[1][1] [4] = 1'b0;
   assign \output_data[1][1] [3] = 1'b0;
   assign \output_data[1][1] [2] = 1'b0;
   assign \output_data[1][1] [1] = 1'b0;
   assign \output_data[1][1] [0] = 1'b0;
   assign \output_data[1][2] [15] = 1'b0;
   assign \output_data[1][2] [14] = 1'b0;
   assign \output_data[1][2] [13] = 1'b0;
   assign \output_data[1][2] [12] = 1'b0;
   assign \output_data[1][2] [11] = 1'b0;
   assign \output_data[1][2] [10] = 1'b0;
   assign \output_data[1][2] [9] = 1'b0;
   assign \output_data[1][2] [8] = 1'b0;
   assign \output_data[1][2] [7] = 1'b0;
   assign \output_data[1][2] [6] = 1'b0;
   assign \output_data[1][2] [5] = 1'b0;
   assign \output_data[1][2] [4] = 1'b0;
   assign \output_data[1][2] [3] = 1'b0;
   assign \output_data[1][2] [2] = 1'b0;
   assign \output_data[1][2] [1] = 1'b0;
   assign \output_data[1][2] [0] = 1'b0;
   assign \output_data[1][3] [15] = 1'b0;
   assign \output_data[1][3] [14] = 1'b0;
   assign \output_data[1][3] [13] = 1'b0;
   assign \output_data[1][3] [12] = 1'b0;
   assign \output_data[1][3] [11] = 1'b0;
   assign \output_data[1][3] [10] = 1'b0;
   assign \output_data[1][3] [9] = 1'b0;
   assign \output_data[1][3] [8] = 1'b0;
   assign \output_data[1][3] [7] = 1'b0;
   assign \output_data[1][3] [6] = 1'b0;
   assign \output_data[1][3] [5] = 1'b0;
   assign \output_data[1][3] [4] = 1'b0;
   assign \output_data[1][3] [3] = 1'b0;
   assign \output_data[1][3] [2] = 1'b0;
   assign \output_data[1][3] [1] = 1'b0;
   assign \output_data[1][3] [0] = 1'b0;
   assign \output_data[1][4] [15] = 1'b0;
   assign \output_data[1][4] [14] = 1'b0;
   assign \output_data[1][4] [13] = 1'b0;
   assign \output_data[1][4] [12] = 1'b0;
   assign \output_data[1][4] [11] = 1'b0;
   assign \output_data[1][4] [10] = 1'b0;
   assign \output_data[1][4] [9] = 1'b0;
   assign \output_data[1][4] [8] = 1'b0;
   assign \output_data[1][4] [7] = 1'b0;
   assign \output_data[1][4] [6] = 1'b0;
   assign \output_data[1][4] [5] = 1'b0;
   assign \output_data[1][4] [4] = 1'b0;
   assign \output_data[1][4] [3] = 1'b0;
   assign \output_data[1][4] [2] = 1'b0;
   assign \output_data[1][4] [1] = 1'b0;
   assign \output_data[1][4] [0] = 1'b0;
   assign \output_data[2][0] [15] = 1'b0;
   assign \output_data[2][0] [14] = 1'b0;
   assign \output_data[2][0] [13] = 1'b0;
   assign \output_data[2][0] [12] = 1'b0;
   assign \output_data[2][0] [11] = 1'b0;
   assign \output_data[2][0] [10] = 1'b0;
   assign \output_data[2][0] [9] = 1'b0;
   assign \output_data[2][0] [8] = 1'b0;
   assign \output_data[2][0] [7] = 1'b0;
   assign \output_data[2][0] [6] = 1'b0;
   assign \output_data[2][0] [5] = 1'b0;
   assign \output_data[2][0] [4] = 1'b0;
   assign \output_data[2][0] [3] = 1'b0;
   assign \output_data[2][0] [2] = 1'b0;
   assign \output_data[2][0] [1] = 1'b0;
   assign \output_data[2][0] [0] = 1'b0;
   assign \output_data[2][1] [15] = 1'b0;
   assign \output_data[2][1] [14] = 1'b0;
   assign \output_data[2][1] [13] = 1'b0;
   assign \output_data[2][1] [12] = 1'b0;
   assign \output_data[2][1] [11] = 1'b0;
   assign \output_data[2][1] [10] = 1'b0;
   assign \output_data[2][1] [9] = 1'b0;
   assign \output_data[2][1] [8] = 1'b0;
   assign \output_data[2][1] [7] = 1'b0;
   assign \output_data[2][1] [6] = 1'b0;
   assign \output_data[2][1] [5] = 1'b0;
   assign \output_data[2][1] [4] = 1'b0;
   assign \output_data[2][1] [3] = 1'b0;
   assign \output_data[2][1] [2] = 1'b0;
   assign \output_data[2][1] [1] = 1'b0;
   assign \output_data[2][1] [0] = 1'b0;
   assign \output_data[2][2] [15] = 1'b0;
   assign \output_data[2][2] [14] = 1'b0;
   assign \output_data[2][2] [13] = 1'b0;
   assign \output_data[2][2] [12] = 1'b0;
   assign \output_data[2][2] [11] = 1'b0;
   assign \output_data[2][2] [10] = 1'b0;
   assign \output_data[2][2] [9] = 1'b0;
   assign \output_data[2][2] [8] = 1'b0;
   assign \output_data[2][2] [7] = 1'b0;
   assign \output_data[2][2] [6] = 1'b0;
   assign \output_data[2][2] [5] = 1'b0;
   assign \output_data[2][2] [4] = 1'b0;
   assign \output_data[2][2] [3] = 1'b0;
   assign \output_data[2][2] [2] = 1'b0;
   assign \output_data[2][2] [1] = 1'b0;
   assign \output_data[2][2] [0] = 1'b0;
   assign \output_data[2][3] [15] = 1'b0;
   assign \output_data[2][3] [14] = 1'b0;
   assign \output_data[2][3] [13] = 1'b0;
   assign \output_data[2][3] [12] = 1'b0;
   assign \output_data[2][3] [11] = 1'b0;
   assign \output_data[2][3] [10] = 1'b0;
   assign \output_data[2][3] [9] = 1'b0;
   assign \output_data[2][3] [8] = 1'b0;
   assign \output_data[2][3] [7] = 1'b0;
   assign \output_data[2][3] [6] = 1'b0;
   assign \output_data[2][3] [5] = 1'b0;
   assign \output_data[2][3] [4] = 1'b0;
   assign \output_data[2][3] [3] = 1'b0;
   assign \output_data[2][3] [2] = 1'b0;
   assign \output_data[2][3] [1] = 1'b0;
   assign \output_data[2][3] [0] = 1'b0;
   assign \output_data[2][4] [15] = 1'b0;
   assign \output_data[2][4] [14] = 1'b0;
   assign \output_data[2][4] [13] = 1'b0;
   assign \output_data[2][4] [12] = 1'b0;
   assign \output_data[2][4] [11] = 1'b0;
   assign \output_data[2][4] [10] = 1'b0;
   assign \output_data[2][4] [9] = 1'b0;
   assign \output_data[2][4] [8] = 1'b0;
   assign \output_data[2][4] [7] = 1'b0;
   assign \output_data[2][4] [6] = 1'b0;
   assign \output_data[2][4] [5] = 1'b0;
   assign \output_data[2][4] [4] = 1'b0;
   assign \output_data[2][4] [3] = 1'b0;
   assign \output_data[2][4] [2] = 1'b0;
   assign \output_data[2][4] [1] = 1'b0;
   assign \output_data[2][4] [0] = 1'b0;
   assign \output_data[3][0] [15] = 1'b0;
   assign \output_data[3][0] [14] = 1'b0;
   assign \output_data[3][0] [13] = 1'b0;
   assign \output_data[3][0] [12] = 1'b0;
   assign \output_data[3][0] [11] = 1'b0;
   assign \output_data[3][0] [10] = 1'b0;
   assign \output_data[3][0] [9] = 1'b0;
   assign \output_data[3][0] [8] = 1'b0;
   assign \output_data[3][0] [7] = 1'b0;
   assign \output_data[3][0] [6] = 1'b0;
   assign \output_data[3][0] [5] = 1'b0;
   assign \output_data[3][0] [4] = 1'b0;
   assign \output_data[3][0] [3] = 1'b0;
   assign \output_data[3][0] [2] = 1'b0;
   assign \output_data[3][0] [1] = 1'b0;
   assign \output_data[3][0] [0] = 1'b0;
   assign \output_data[3][1] [15] = 1'b0;
   assign \output_data[3][1] [14] = 1'b0;
   assign \output_data[3][1] [13] = 1'b0;
   assign \output_data[3][1] [12] = 1'b0;
   assign \output_data[3][1] [11] = 1'b0;
   assign \output_data[3][1] [10] = 1'b0;
   assign \output_data[3][1] [9] = 1'b0;
   assign \output_data[3][1] [8] = 1'b0;
   assign \output_data[3][1] [7] = 1'b0;
   assign \output_data[3][1] [6] = 1'b0;
   assign \output_data[3][1] [5] = 1'b0;
   assign \output_data[3][1] [4] = 1'b0;
   assign \output_data[3][1] [3] = 1'b0;
   assign \output_data[3][1] [2] = 1'b0;
   assign \output_data[3][1] [1] = 1'b0;
   assign \output_data[3][1] [0] = 1'b0;
   assign \output_data[3][2] [15] = 1'b0;
   assign \output_data[3][2] [14] = 1'b0;
   assign \output_data[3][2] [13] = 1'b0;
   assign \output_data[3][2] [12] = 1'b0;
   assign \output_data[3][2] [11] = 1'b0;
   assign \output_data[3][2] [10] = 1'b0;
   assign \output_data[3][2] [9] = 1'b0;
   assign \output_data[3][2] [8] = 1'b0;
   assign \output_data[3][2] [7] = 1'b0;
   assign \output_data[3][2] [6] = 1'b0;
   assign \output_data[3][2] [5] = 1'b0;
   assign \output_data[3][2] [4] = 1'b0;
   assign \output_data[3][2] [3] = 1'b0;
   assign \output_data[3][2] [2] = 1'b0;
   assign \output_data[3][2] [1] = 1'b0;
   assign \output_data[3][2] [0] = 1'b0;
   assign \output_data[3][3] [15] = 1'b0;
   assign \output_data[3][3] [14] = 1'b0;
   assign \output_data[3][3] [13] = 1'b0;
   assign \output_data[3][3] [12] = 1'b0;
   assign \output_data[3][3] [11] = 1'b0;
   assign \output_data[3][3] [10] = 1'b0;
   assign \output_data[3][3] [9] = 1'b0;
   assign \output_data[3][3] [8] = 1'b0;
   assign \output_data[3][3] [7] = 1'b0;
   assign \output_data[3][3] [6] = 1'b0;
   assign \output_data[3][3] [5] = 1'b0;
   assign \output_data[3][3] [4] = 1'b0;
   assign \output_data[3][3] [3] = 1'b0;
   assign \output_data[3][3] [2] = 1'b0;
   assign \output_data[3][3] [1] = 1'b0;
   assign \output_data[3][3] [0] = 1'b0;
   assign \output_data[3][4] [15] = 1'b0;
   assign \output_data[3][4] [14] = 1'b0;
   assign \output_data[3][4] [13] = 1'b0;
   assign \output_data[3][4] [12] = 1'b0;
   assign \output_data[3][4] [11] = 1'b0;
   assign \output_data[3][4] [10] = 1'b0;
   assign \output_data[3][4] [9] = 1'b0;
   assign \output_data[3][4] [8] = 1'b0;
   assign \output_data[3][4] [7] = 1'b0;
   assign \output_data[3][4] [6] = 1'b0;
   assign \output_data[3][4] [5] = 1'b0;
   assign \output_data[3][4] [4] = 1'b0;
   assign \output_data[3][4] [3] = 1'b0;
   assign \output_data[3][4] [2] = 1'b0;
   assign \output_data[3][4] [1] = 1'b0;
   assign \output_data[3][4] [0] = 1'b0;
   assign \output_data[4][0] [15] = 1'b0;
   assign \output_data[4][0] [14] = 1'b0;
   assign \output_data[4][0] [13] = 1'b0;
   assign \output_data[4][0] [12] = 1'b0;
   assign \output_data[4][0] [11] = 1'b0;
   assign \output_data[4][0] [10] = 1'b0;
   assign \output_data[4][0] [9] = 1'b0;
   assign \output_data[4][0] [8] = 1'b0;
   assign \output_data[4][0] [7] = 1'b0;
   assign \output_data[4][0] [6] = 1'b0;
   assign \output_data[4][0] [5] = 1'b0;
   assign \output_data[4][0] [4] = 1'b0;
   assign \output_data[4][0] [3] = 1'b0;
   assign \output_data[4][0] [2] = 1'b0;
   assign \output_data[4][0] [1] = 1'b0;
   assign \output_data[4][0] [0] = 1'b0;
   assign \output_data[4][1] [15] = 1'b0;
   assign \output_data[4][1] [14] = 1'b0;
   assign \output_data[4][1] [13] = 1'b0;
   assign \output_data[4][1] [12] = 1'b0;
   assign \output_data[4][1] [11] = 1'b0;
   assign \output_data[4][1] [10] = 1'b0;
   assign \output_data[4][1] [9] = 1'b0;
   assign \output_data[4][1] [8] = 1'b0;
   assign \output_data[4][1] [7] = 1'b0;
   assign \output_data[4][1] [6] = 1'b0;
   assign \output_data[4][1] [5] = 1'b0;
   assign \output_data[4][1] [4] = 1'b0;
   assign \output_data[4][1] [3] = 1'b0;
   assign \output_data[4][1] [2] = 1'b0;
   assign \output_data[4][1] [1] = 1'b0;
   assign \output_data[4][1] [0] = 1'b0;
   assign \output_data[4][2] [15] = 1'b0;
   assign \output_data[4][2] [14] = 1'b0;
   assign \output_data[4][2] [13] = 1'b0;
   assign \output_data[4][2] [12] = 1'b0;
   assign \output_data[4][2] [11] = 1'b0;
   assign \output_data[4][2] [10] = 1'b0;
   assign \output_data[4][2] [9] = 1'b0;
   assign \output_data[4][2] [8] = 1'b0;
   assign \output_data[4][2] [7] = 1'b0;
   assign \output_data[4][2] [6] = 1'b0;
   assign \output_data[4][2] [5] = 1'b0;
   assign \output_data[4][2] [4] = 1'b0;
   assign \output_data[4][2] [3] = 1'b0;
   assign \output_data[4][2] [2] = 1'b0;
   assign \output_data[4][2] [1] = 1'b0;
   assign \output_data[4][2] [0] = 1'b0;
   assign \output_data[4][3] [15] = 1'b0;
   assign \output_data[4][3] [14] = 1'b0;
   assign \output_data[4][3] [13] = 1'b0;
   assign \output_data[4][3] [12] = 1'b0;
   assign \output_data[4][3] [11] = 1'b0;
   assign \output_data[4][3] [10] = 1'b0;
   assign \output_data[4][3] [9] = 1'b0;
   assign \output_data[4][3] [8] = 1'b0;
   assign \output_data[4][3] [7] = 1'b0;
   assign \output_data[4][3] [6] = 1'b0;
   assign \output_data[4][3] [5] = 1'b0;
   assign \output_data[4][3] [4] = 1'b0;
   assign \output_data[4][3] [3] = 1'b0;
   assign \output_data[4][3] [2] = 1'b0;
   assign \output_data[4][3] [1] = 1'b0;
   assign \output_data[4][3] [0] = 1'b0;
   assign \output_data[4][4] [15] = 1'b0;
   assign \output_data[4][4] [14] = 1'b0;
   assign \output_data[4][4] [13] = 1'b0;
   assign \output_data[4][4] [12] = 1'b0;
   assign \output_data[4][4] [11] = 1'b0;
   assign \output_data[4][4] [10] = 1'b0;
   assign \output_data[4][4] [9] = 1'b0;
   assign \output_data[4][4] [8] = 1'b0;
   assign \output_data[4][4] [7] = 1'b0;
   assign \output_data[4][4] [6] = 1'b0;
   assign \output_data[4][4] [5] = 1'b0;
   assign \output_data[4][4] [4] = 1'b0;
   assign \output_data[4][4] [3] = 1'b0;
   assign \output_data[4][4] [2] = 1'b0;
   assign \output_data[4][4] [1] = 1'b0;
   assign \output_data[4][4] [0] = 1'b0;
   assign finish = 1'b0;

   DFF_X1 finish_flag_reg__0 (.D(1'b0), .CK(n_27_0), .Q(1'b0), .QN());
   INV_X1 i_27_0_0 (.A(clk), .ZN(n_27_0));
endmodule

module datapath__0_73(p_0, p_1, inner_address);
   input [5:0]p_0;
   input [15:0]p_1;
   output [15:0]inner_address;

   HA_X1 i_2 (.A(p_0[0]), .B(p_1[5]), .CO(n_3), .S(n_2));
   HA_X1 i_3 (.A(p_1[6]), .B(n_3), .CO(n_5), .S(n_4));
   HA_X1 i_4 (.A(p_1[7]), .B(n_5), .CO(n_7), .S(n_6));
   HA_X1 i_5 (.A(p_1[8]), .B(n_1), .CO(n_9), .S(n_8));
   HA_X1 i_6 (.A(p_1[9]), .B(n_1), .CO(n_11), .S(n_10));
   HA_X1 i_7 (.A(p_1[10]), .B(n_1), .CO(n_13), .S(n_12));
   HA_X1 i_8 (.A(p_1[11]), .B(n_1), .CO(n_15), .S(n_14));
   HA_X1 i_9 (.A(p_1[12]), .B(n_1), .CO(n_17), .S(n_16));
   HA_X1 i_10 (.A(p_1[13]), .B(n_1), .CO(n_19), .S(n_18));
   HA_X1 i_11 (.A(p_1[14]), .B(n_1), .CO(n_21), .S(n_20));
   HA_X1 i_14 (.A(p_0[0]), .B(p_1[0]), .CO(n_24), .S(inner_address[0]));
   HA_X1 i_15 (.A(p_1[1]), .B(n_24), .CO(n_25), .S(inner_address[1]));
   HA_X1 i_16 (.A(p_1[2]), .B(n_25), .CO(n_26), .S(inner_address[2]));
   FA_X1 i_17 (.A(p_1[3]), .B(p_0[0]), .CI(n_26), .CO(n_27), .S(inner_address[3]));
   FA_X1 i_18 (.A(n_0), .B(n_1), .CI(n_27), .CO(n_28), .S(inner_address[4]));
   FA_X1 i_19 (.A(n_2), .B(n_1), .CI(n_28), .CO(n_29), .S(inner_address[5]));
   FA_X1 i_20 (.A(n_1), .B(n_4), .CI(n_29), .CO(n_30), .S(inner_address[6]));
   FA_X1 i_21 (.A(n_1), .B(n_6), .CI(n_30), .CO(n_31), .S(inner_address[7]));
   FA_X1 i_22 (.A(n_7), .B(n_8), .CI(n_31), .CO(n_32), .S(inner_address[8]));
   FA_X1 i_23 (.A(n_9), .B(n_10), .CI(n_32), .CO(n_33), .S(inner_address[9]));
   FA_X1 i_24 (.A(n_11), .B(n_12), .CI(n_33), .CO(n_34), .S(inner_address[10]));
   FA_X1 i_25 (.A(n_13), .B(n_14), .CI(n_34), .CO(n_35), .S(inner_address[11]));
   FA_X1 i_26 (.A(n_15), .B(n_16), .CI(n_35), .CO(n_36), .S(inner_address[12]));
   FA_X1 i_27 (.A(n_17), .B(n_18), .CI(n_36), .CO(n_37), .S(inner_address[13]));
   FA_X1 i_28 (.A(n_19), .B(n_20), .CI(n_37), .CO(n_38), .S(inner_address[14]));
   XNOR2_X1 i_0 (.A(n_23), .B(n_22), .ZN(inner_address[15]));
   XNOR2_X1 i_1 (.A(n_21), .B(n_38), .ZN(n_22));
   XNOR2_X1 i_12 (.A(p_1[15]), .B(p_1[4]), .ZN(n_23));
   INV_X1 i_13 (.A(p_1[4]), .ZN(n_1));
   INV_X1 i_29 (.A(p_0[0]), .ZN(n_0));
endmodule

module DMA(start, reset, finish_read, clk, address, offset, 
      read_write_filter_bias, filter_number, \CNN_output_data[0][0] , 
      \CNN_output_data[0][1] , \CNN_output_data[0][2] , \CNN_output_data[0][3] , 
      \CNN_output_data[0][4] , \CNN_output_data[1][0] , \CNN_output_data[1][1] , 
      \CNN_output_data[1][2] , \CNN_output_data[1][3] , \CNN_output_data[1][4] , 
      \CNN_output_data[2][0] , \CNN_output_data[2][1] , \CNN_output_data[2][2] , 
      \CNN_output_data[2][3] , \CNN_output_data[2][4] , \CNN_output_data[3][0] , 
      \CNN_output_data[3][1] , \CNN_output_data[3][2] , \CNN_output_data[3][3] , 
      \CNN_output_data[3][4] , \CNN_output_data[4][0] , \CNN_output_data[4][1] , 
      \CNN_output_data[4][2] , \CNN_output_data[4][3] , \CNN_output_data[4][4] , 
      CNN_input_data, RAM_address, RAM_offset, RAM_write, RAM_output_data, 
      \RAM_input_data[0][0] , \RAM_input_data[0][1] , \RAM_input_data[0][2] , 
      \RAM_input_data[0][3] , \RAM_input_data[0][4] , \RAM_input_data[1][0] , 
      \RAM_input_data[1][1] , \RAM_input_data[1][2] , \RAM_input_data[1][3] , 
      \RAM_input_data[1][4] , \RAM_input_data[2][0] , \RAM_input_data[2][1] , 
      \RAM_input_data[2][2] , \RAM_input_data[2][3] , \RAM_input_data[2][4] , 
      \RAM_input_data[3][0] , \RAM_input_data[3][1] , \RAM_input_data[3][2] , 
      \RAM_input_data[3][3] , \RAM_input_data[3][4] , \RAM_input_data[4][0] , 
      \RAM_input_data[4][1] , \RAM_input_data[4][2] , \RAM_input_data[4][3] , 
      \RAM_input_data[4][4] , RAM_finish, RAM_enable, FB_write, 
      \FB_filter[0][0] , \FB_filter[0][1] , \FB_filter[0][2] , \FB_filter[0][3] , 
      \FB_filter[0][4] , \FB_filter[1][0] , \FB_filter[1][1] , \FB_filter[1][2] , 
      \FB_filter[1][3] , \FB_filter[1][4] , \FB_filter[2][0] , \FB_filter[2][1] , 
      \FB_filter[2][2] , \FB_filter[2][3] , \FB_filter[2][4] , \FB_filter[3][0] , 
      \FB_filter[3][1] , \FB_filter[3][2] , \FB_filter[3][3] , \FB_filter[3][4] , 
      \FB_filter[4][0] , \FB_filter[4][1] , \FB_filter[4][2] , \FB_filter[4][3] , 
      \FB_filter[4][4] , FB_index_filter, \FB_bias[0] , \FB_bias[1] , 
      \FB_bias[2] , \FB_bias[3] , \FB_bias[4] , \FB_bias[5] , \FB_bias[6] , 
      \FB_bias[7] , \FB_bias[8] , \FB_bias[9] , \FB_bias[10] , \FB_bias[11] , 
      \FB_bias[12] , \FB_bias[13] , \FB_bias[14] , \FB_bias[15] , \FB_bias[16] , 
      \FB_bias[17] , \FB_bias[18] , \FB_bias[19] , \FB_bias[20] , \FB_bias[21] , 
      \FB_bias[22] , \FB_bias[23] , \FB_bias[24] , \FB_bias[25] , \FB_bias[26] , 
      \FB_bias[27] , \FB_bias[28] , \FB_bias[29] , \FB_bias[30] , \FB_bias[31] , 
      \FB_bias[32] , \FB_bias[33] , \FB_bias[34] , \FB_bias[35] , \FB_bias[36] , 
      \FB_bias[37] , \FB_bias[38] , \FB_bias[39] , \FB_bias[40] , \FB_bias[41] , 
      \FB_bias[42] , \FB_bias[43] , \FB_bias[44] , \FB_bias[45] , \FB_bias[46] , 
      \FB_bias[47] , \FB_bias[48] , \FB_bias[49] , \FB_bias[50] , \FB_bias[51] , 
      \FB_bias[52] , \FB_bias[53] , \FB_bias[54] , \FB_bias[55] , \FB_bias[56] , 
      \FB_bias[57] , \FB_bias[58] , \FB_bias[59] , \FB_bias[60] , \FB_bias[61] , 
      \FB_bias[62] , \FB_bias[63] , \FB_bias[64] , \FB_bias[65] , \FB_bias[66] , 
      \FB_bias[67] , \FB_bias[68] , \FB_bias[69] , \FB_bias[70] , \FB_bias[71] , 
      \FB_bias[72] , \FB_bias[73] , \FB_bias[74] , \FB_bias[75] , \FB_bias[76] , 
      \FB_bias[77] , \FB_bias[78] , \FB_bias[79] , \FB_bias[80] , \FB_bias[81] , 
      \FB_bias[82] , \FB_bias[83] , \FB_bias[84] , \FB_bias[85] , \FB_bias[86] , 
      \FB_bias[87] , \FB_bias[88] , \FB_bias[89] , \FB_bias[90] , \FB_bias[91] , 
      \FB_bias[92] , \FB_bias[93] , \FB_bias[94] , \FB_bias[95] , \FB_bias[96] , 
      \FB_bias[97] , \FB_bias[98] , \FB_bias[99] , \FB_bias[100] , 
      \FB_bias[101] , \FB_bias[102] , \FB_bias[103] , \FB_bias[104] , 
      \FB_bias[105] , \FB_bias[106] , \FB_bias[107] , \FB_bias[108] , 
      \FB_bias[109] , \FB_bias[110] , \FB_bias[111] , \FB_bias[112] , 
      \FB_bias[113] , \FB_bias[114] , \FB_bias[115] , \FB_bias[116] , 
      \FB_bias[117] , \FB_bias[118] , \FB_bias[119] , FB_bias_or_filter);
   input start;
   input reset;
   output finish_read;
   input clk;
   input [15:0]address;
   input [15:0]offset;
   input [1:0]read_write_filter_bias;
   input [15:0]filter_number;
   output [15:0]\CNN_output_data[0][0] ;
   output [15:0]\CNN_output_data[0][1] ;
   output [15:0]\CNN_output_data[0][2] ;
   output [15:0]\CNN_output_data[0][3] ;
   output [15:0]\CNN_output_data[0][4] ;
   output [15:0]\CNN_output_data[1][0] ;
   output [15:0]\CNN_output_data[1][1] ;
   output [15:0]\CNN_output_data[1][2] ;
   output [15:0]\CNN_output_data[1][3] ;
   output [15:0]\CNN_output_data[1][4] ;
   output [15:0]\CNN_output_data[2][0] ;
   output [15:0]\CNN_output_data[2][1] ;
   output [15:0]\CNN_output_data[2][2] ;
   output [15:0]\CNN_output_data[2][3] ;
   output [15:0]\CNN_output_data[2][4] ;
   output [15:0]\CNN_output_data[3][0] ;
   output [15:0]\CNN_output_data[3][1] ;
   output [15:0]\CNN_output_data[3][2] ;
   output [15:0]\CNN_output_data[3][3] ;
   output [15:0]\CNN_output_data[3][4] ;
   output [15:0]\CNN_output_data[4][0] ;
   output [15:0]\CNN_output_data[4][1] ;
   output [15:0]\CNN_output_data[4][2] ;
   output [15:0]\CNN_output_data[4][3] ;
   output [15:0]\CNN_output_data[4][4] ;
   input [15:0]CNN_input_data;
   output [15:0]RAM_address;
   output [15:0]RAM_offset;
   output RAM_write;
   output [15:0]RAM_output_data;
   input [15:0]\RAM_input_data[0][0] ;
   input [15:0]\RAM_input_data[0][1] ;
   input [15:0]\RAM_input_data[0][2] ;
   input [15:0]\RAM_input_data[0][3] ;
   input [15:0]\RAM_input_data[0][4] ;
   input [15:0]\RAM_input_data[1][0] ;
   input [15:0]\RAM_input_data[1][1] ;
   input [15:0]\RAM_input_data[1][2] ;
   input [15:0]\RAM_input_data[1][3] ;
   input [15:0]\RAM_input_data[1][4] ;
   input [15:0]\RAM_input_data[2][0] ;
   input [15:0]\RAM_input_data[2][1] ;
   input [15:0]\RAM_input_data[2][2] ;
   input [15:0]\RAM_input_data[2][3] ;
   input [15:0]\RAM_input_data[2][4] ;
   input [15:0]\RAM_input_data[3][0] ;
   input [15:0]\RAM_input_data[3][1] ;
   input [15:0]\RAM_input_data[3][2] ;
   input [15:0]\RAM_input_data[3][3] ;
   input [15:0]\RAM_input_data[3][4] ;
   input [15:0]\RAM_input_data[4][0] ;
   input [15:0]\RAM_input_data[4][1] ;
   input [15:0]\RAM_input_data[4][2] ;
   input [15:0]\RAM_input_data[4][3] ;
   input [15:0]\RAM_input_data[4][4] ;
   input RAM_finish;
   output RAM_enable;
   output FB_write;
   output [15:0]\FB_filter[0][0] ;
   output [15:0]\FB_filter[0][1] ;
   output [15:0]\FB_filter[0][2] ;
   output [15:0]\FB_filter[0][3] ;
   output [15:0]\FB_filter[0][4] ;
   output [15:0]\FB_filter[1][0] ;
   output [15:0]\FB_filter[1][1] ;
   output [15:0]\FB_filter[1][2] ;
   output [15:0]\FB_filter[1][3] ;
   output [15:0]\FB_filter[1][4] ;
   output [15:0]\FB_filter[2][0] ;
   output [15:0]\FB_filter[2][1] ;
   output [15:0]\FB_filter[2][2] ;
   output [15:0]\FB_filter[2][3] ;
   output [15:0]\FB_filter[2][4] ;
   output [15:0]\FB_filter[3][0] ;
   output [15:0]\FB_filter[3][1] ;
   output [15:0]\FB_filter[3][2] ;
   output [15:0]\FB_filter[3][3] ;
   output [15:0]\FB_filter[3][4] ;
   output [15:0]\FB_filter[4][0] ;
   output [15:0]\FB_filter[4][1] ;
   output [15:0]\FB_filter[4][2] ;
   output [15:0]\FB_filter[4][3] ;
   output [15:0]\FB_filter[4][4] ;
   output [15:0]FB_index_filter;
   output [15:0]\FB_bias[0] ;
   output [15:0]\FB_bias[1] ;
   output [15:0]\FB_bias[2] ;
   output [15:0]\FB_bias[3] ;
   output [15:0]\FB_bias[4] ;
   output [15:0]\FB_bias[5] ;
   output [15:0]\FB_bias[6] ;
   output [15:0]\FB_bias[7] ;
   output [15:0]\FB_bias[8] ;
   output [15:0]\FB_bias[9] ;
   output [15:0]\FB_bias[10] ;
   output [15:0]\FB_bias[11] ;
   output [15:0]\FB_bias[12] ;
   output [15:0]\FB_bias[13] ;
   output [15:0]\FB_bias[14] ;
   output [15:0]\FB_bias[15] ;
   output [15:0]\FB_bias[16] ;
   output [15:0]\FB_bias[17] ;
   output [15:0]\FB_bias[18] ;
   output [15:0]\FB_bias[19] ;
   output [15:0]\FB_bias[20] ;
   output [15:0]\FB_bias[21] ;
   output [15:0]\FB_bias[22] ;
   output [15:0]\FB_bias[23] ;
   output [15:0]\FB_bias[24] ;
   output [15:0]\FB_bias[25] ;
   output [15:0]\FB_bias[26] ;
   output [15:0]\FB_bias[27] ;
   output [15:0]\FB_bias[28] ;
   output [15:0]\FB_bias[29] ;
   output [15:0]\FB_bias[30] ;
   output [15:0]\FB_bias[31] ;
   output [15:0]\FB_bias[32] ;
   output [15:0]\FB_bias[33] ;
   output [15:0]\FB_bias[34] ;
   output [15:0]\FB_bias[35] ;
   output [15:0]\FB_bias[36] ;
   output [15:0]\FB_bias[37] ;
   output [15:0]\FB_bias[38] ;
   output [15:0]\FB_bias[39] ;
   output [15:0]\FB_bias[40] ;
   output [15:0]\FB_bias[41] ;
   output [15:0]\FB_bias[42] ;
   output [15:0]\FB_bias[43] ;
   output [15:0]\FB_bias[44] ;
   output [15:0]\FB_bias[45] ;
   output [15:0]\FB_bias[46] ;
   output [15:0]\FB_bias[47] ;
   output [15:0]\FB_bias[48] ;
   output [15:0]\FB_bias[49] ;
   output [15:0]\FB_bias[50] ;
   output [15:0]\FB_bias[51] ;
   output [15:0]\FB_bias[52] ;
   output [15:0]\FB_bias[53] ;
   output [15:0]\FB_bias[54] ;
   output [15:0]\FB_bias[55] ;
   output [15:0]\FB_bias[56] ;
   output [15:0]\FB_bias[57] ;
   output [15:0]\FB_bias[58] ;
   output [15:0]\FB_bias[59] ;
   output [15:0]\FB_bias[60] ;
   output [15:0]\FB_bias[61] ;
   output [15:0]\FB_bias[62] ;
   output [15:0]\FB_bias[63] ;
   output [15:0]\FB_bias[64] ;
   output [15:0]\FB_bias[65] ;
   output [15:0]\FB_bias[66] ;
   output [15:0]\FB_bias[67] ;
   output [15:0]\FB_bias[68] ;
   output [15:0]\FB_bias[69] ;
   output [15:0]\FB_bias[70] ;
   output [15:0]\FB_bias[71] ;
   output [15:0]\FB_bias[72] ;
   output [15:0]\FB_bias[73] ;
   output [15:0]\FB_bias[74] ;
   output [15:0]\FB_bias[75] ;
   output [15:0]\FB_bias[76] ;
   output [15:0]\FB_bias[77] ;
   output [15:0]\FB_bias[78] ;
   output [15:0]\FB_bias[79] ;
   output [15:0]\FB_bias[80] ;
   output [15:0]\FB_bias[81] ;
   output [15:0]\FB_bias[82] ;
   output [15:0]\FB_bias[83] ;
   output [15:0]\FB_bias[84] ;
   output [15:0]\FB_bias[85] ;
   output [15:0]\FB_bias[86] ;
   output [15:0]\FB_bias[87] ;
   output [15:0]\FB_bias[88] ;
   output [15:0]\FB_bias[89] ;
   output [15:0]\FB_bias[90] ;
   output [15:0]\FB_bias[91] ;
   output [15:0]\FB_bias[92] ;
   output [15:0]\FB_bias[93] ;
   output [15:0]\FB_bias[94] ;
   output [15:0]\FB_bias[95] ;
   output [15:0]\FB_bias[96] ;
   output [15:0]\FB_bias[97] ;
   output [15:0]\FB_bias[98] ;
   output [15:0]\FB_bias[99] ;
   output [15:0]\FB_bias[100] ;
   output [15:0]\FB_bias[101] ;
   output [15:0]\FB_bias[102] ;
   output [15:0]\FB_bias[103] ;
   output [15:0]\FB_bias[104] ;
   output [15:0]\FB_bias[105] ;
   output [15:0]\FB_bias[106] ;
   output [15:0]\FB_bias[107] ;
   output [15:0]\FB_bias[108] ;
   output [15:0]\FB_bias[109] ;
   output [15:0]\FB_bias[110] ;
   output [15:0]\FB_bias[111] ;
   output [15:0]\FB_bias[112] ;
   output [15:0]\FB_bias[113] ;
   output [15:0]\FB_bias[114] ;
   output [15:0]\FB_bias[115] ;
   output [15:0]\FB_bias[116] ;
   output [15:0]\FB_bias[117] ;
   output [15:0]\FB_bias[118] ;
   output [15:0]\FB_bias[119] ;
   output FB_bias_or_filter;

   wire n_1_29;
   wire n_1_30;
   wire n_1_31;
   wire n_1_32;
   wire n_1_33;
   wire n_1_34;
   wire n_1_35;
   wire n_1_36;
   wire n_1_37;
   wire n_1_38;
   wire n_1_39;
   wire n_1_40;
   wire n_1_41;
   wire n_1_42;
   wire n_1_43;
   wire n_1_44;
   wire n_1_0_1;
   wire n_1_0_4;
   wire n_1_0_0;
   wire n_1_0_5;
   wire n_1_0_2;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_0_6;
   wire n_1_4;
   wire n_1_5;
   wire n_1_77;
   wire n_1_0_7;
   wire n_1_6;
   wire n_1_0_8;
   wire n_1_7;
   wire n_1_0_9;
   wire n_1_8;
   wire n_1_0_10;
   wire n_1_9;
   wire n_1_0_11;
   wire n_1_10;
   wire n_1_0_12;
   wire n_1_11;
   wire n_1_0_13;
   wire n_1_12;
   wire n_1_0_14;
   wire n_1_13;
   wire n_1_0_15;
   wire n_1_14;
   wire n_1_0_16;
   wire n_1_15;
   wire n_1_0_17;
   wire n_1_16;
   wire n_1_0_18;
   wire n_1_17;
   wire n_1_0_19;
   wire n_1_18;
   wire n_1_0_20;
   wire n_1_19;
   wire n_1_0_21;
   wire n_1_20;
   wire n_1_0_22;
   wire n_1_0_23;
   wire n_1_0_24;
   wire n_1_0_25;
   wire n_1_61;
   wire n_1_0_26;
   wire n_1_62;
   wire n_1_0_27;
   wire n_1_63;
   wire n_1_0_28;
   wire n_1_64;
   wire n_1_0_29;
   wire n_1_65;
   wire n_1_0_30;
   wire n_1_66;
   wire n_1_0_31;
   wire n_1_67;
   wire n_1_0_32;
   wire n_1_68;
   wire n_1_0_33;
   wire n_1_69;
   wire n_1_0_34;
   wire n_1_70;
   wire n_1_0_35;
   wire n_1_71;
   wire n_1_0_36;
   wire n_1_72;
   wire n_1_0_37;
   wire n_1_73;
   wire n_1_0_38;
   wire n_1_74;
   wire n_1_0_39;
   wire n_1_75;
   wire n_1_0_40;
   wire n_1_76;
   wire n_1_0_41;
   wire n_1_21;
   wire n_1_22;
   wire n_1_23;
   wire n_1_24;
   wire n_1_25;
   wire n_1_26;
   wire n_1_27;
   wire n_1_28;
   wire n_1_45;
   wire n_1_46;
   wire n_1_47;
   wire n_1_48;
   wire n_1_49;
   wire n_1_50;
   wire n_1_51;
   wire n_1_52;
   wire n_1_0_42;
   wire n_1_0_3;
   wire n_1_54;
   wire n_1_53;
   wire n_1_0_43;
   wire n_1_0_44;
   wire n_1_0_45;
   wire n_1_78;
   wire n_1_0_46;
   wire n_1_0_47;
   wire n_1_0_48;
   wire n_1_55;
   wire n_1_0_49;
   wire n_1_0_50;
   wire n_1_0_51;
   wire n_1_0_52;
   wire n_1_0_53;
   wire n_1_0_54;
   wire n_1_56;
   wire n_1_57;
   wire [31:0]biasCounter;
   wire n_1_58;
   wire [15:0]inner_address;
   wire n_1_59;
   wire n_1_60;
   wire n_0_0;
   wire n_0_1_0;
   wire n_0_1_1;
   wire n_0_16;
   wire n_0_15;
   wire n_0_14;
   wire n_0_13;
   wire n_0_12;
   wire n_0_11;
   wire n_0_10;
   wire n_0_9;
   wire n_0_8;
   wire n_0_7;
   wire n_0_6;
   wire n_0_5;
   wire n_0_4;
   wire n_0_3;
   wire n_0_2;
   wire n_0_1;

   assign \FB_filter[0][0] [15] = 1'b0;
   assign \FB_filter[0][0] [14] = 1'b0;
   assign \FB_filter[0][0] [13] = 1'b0;
   assign \FB_filter[0][0] [12] = 1'b0;
   assign \FB_filter[0][0] [11] = 1'b0;
   assign \FB_filter[0][0] [10] = 1'b0;
   assign \FB_filter[0][0] [9] = 1'b0;
   assign \FB_filter[0][0] [8] = 1'b0;
   assign \FB_filter[0][0] [7] = 1'b0;
   assign \FB_filter[0][0] [6] = 1'b0;
   assign \FB_filter[0][0] [5] = 1'b0;
   assign \FB_filter[0][0] [4] = 1'b0;
   assign \FB_filter[0][0] [3] = 1'b0;
   assign \FB_filter[0][0] [2] = 1'b0;
   assign \FB_filter[0][0] [1] = 1'b0;
   assign \FB_filter[0][0] [0] = 1'b0;
   assign \FB_filter[0][1] [15] = 1'b0;
   assign \FB_filter[0][1] [14] = 1'b0;
   assign \FB_filter[0][1] [13] = 1'b0;
   assign \FB_filter[0][1] [12] = 1'b0;
   assign \FB_filter[0][1] [11] = 1'b0;
   assign \FB_filter[0][1] [10] = 1'b0;
   assign \FB_filter[0][1] [9] = 1'b0;
   assign \FB_filter[0][1] [8] = 1'b0;
   assign \FB_filter[0][1] [7] = 1'b0;
   assign \FB_filter[0][1] [6] = 1'b0;
   assign \FB_filter[0][1] [5] = 1'b0;
   assign \FB_filter[0][1] [4] = 1'b0;
   assign \FB_filter[0][1] [3] = 1'b0;
   assign \FB_filter[0][1] [2] = 1'b0;
   assign \FB_filter[0][1] [1] = 1'b0;
   assign \FB_filter[0][1] [0] = 1'b0;
   assign \FB_filter[0][2] [15] = 1'b0;
   assign \FB_filter[0][2] [14] = 1'b0;
   assign \FB_filter[0][2] [13] = 1'b0;
   assign \FB_filter[0][2] [12] = 1'b0;
   assign \FB_filter[0][2] [11] = 1'b0;
   assign \FB_filter[0][2] [10] = 1'b0;
   assign \FB_filter[0][2] [9] = 1'b0;
   assign \FB_filter[0][2] [8] = 1'b0;
   assign \FB_filter[0][2] [7] = 1'b0;
   assign \FB_filter[0][2] [6] = 1'b0;
   assign \FB_filter[0][2] [5] = 1'b0;
   assign \FB_filter[0][2] [4] = 1'b0;
   assign \FB_filter[0][2] [3] = 1'b0;
   assign \FB_filter[0][2] [2] = 1'b0;
   assign \FB_filter[0][2] [1] = 1'b0;
   assign \FB_filter[0][2] [0] = 1'b0;
   assign \FB_filter[0][3] [15] = 1'b0;
   assign \FB_filter[0][3] [14] = 1'b0;
   assign \FB_filter[0][3] [13] = 1'b0;
   assign \FB_filter[0][3] [12] = 1'b0;
   assign \FB_filter[0][3] [11] = 1'b0;
   assign \FB_filter[0][3] [10] = 1'b0;
   assign \FB_filter[0][3] [9] = 1'b0;
   assign \FB_filter[0][3] [8] = 1'b0;
   assign \FB_filter[0][3] [7] = 1'b0;
   assign \FB_filter[0][3] [6] = 1'b0;
   assign \FB_filter[0][3] [5] = 1'b0;
   assign \FB_filter[0][3] [4] = 1'b0;
   assign \FB_filter[0][3] [3] = 1'b0;
   assign \FB_filter[0][3] [2] = 1'b0;
   assign \FB_filter[0][3] [1] = 1'b0;
   assign \FB_filter[0][3] [0] = 1'b0;
   assign \FB_filter[0][4] [15] = 1'b0;
   assign \FB_filter[0][4] [14] = 1'b0;
   assign \FB_filter[0][4] [13] = 1'b0;
   assign \FB_filter[0][4] [12] = 1'b0;
   assign \FB_filter[0][4] [11] = 1'b0;
   assign \FB_filter[0][4] [10] = 1'b0;
   assign \FB_filter[0][4] [9] = 1'b0;
   assign \FB_filter[0][4] [8] = 1'b0;
   assign \FB_filter[0][4] [7] = 1'b0;
   assign \FB_filter[0][4] [6] = 1'b0;
   assign \FB_filter[0][4] [5] = 1'b0;
   assign \FB_filter[0][4] [4] = 1'b0;
   assign \FB_filter[0][4] [3] = 1'b0;
   assign \FB_filter[0][4] [2] = 1'b0;
   assign \FB_filter[0][4] [1] = 1'b0;
   assign \FB_filter[0][4] [0] = 1'b0;
   assign \FB_filter[1][0] [15] = 1'b0;
   assign \FB_filter[1][0] [14] = 1'b0;
   assign \FB_filter[1][0] [13] = 1'b0;
   assign \FB_filter[1][0] [12] = 1'b0;
   assign \FB_filter[1][0] [11] = 1'b0;
   assign \FB_filter[1][0] [10] = 1'b0;
   assign \FB_filter[1][0] [9] = 1'b0;
   assign \FB_filter[1][0] [8] = 1'b0;
   assign \FB_filter[1][0] [7] = 1'b0;
   assign \FB_filter[1][0] [6] = 1'b0;
   assign \FB_filter[1][0] [5] = 1'b0;
   assign \FB_filter[1][0] [4] = 1'b0;
   assign \FB_filter[1][0] [3] = 1'b0;
   assign \FB_filter[1][0] [2] = 1'b0;
   assign \FB_filter[1][0] [1] = 1'b0;
   assign \FB_filter[1][0] [0] = 1'b0;
   assign \FB_filter[1][1] [15] = 1'b0;
   assign \FB_filter[1][1] [14] = 1'b0;
   assign \FB_filter[1][1] [13] = 1'b0;
   assign \FB_filter[1][1] [12] = 1'b0;
   assign \FB_filter[1][1] [11] = 1'b0;
   assign \FB_filter[1][1] [10] = 1'b0;
   assign \FB_filter[1][1] [9] = 1'b0;
   assign \FB_filter[1][1] [8] = 1'b0;
   assign \FB_filter[1][1] [7] = 1'b0;
   assign \FB_filter[1][1] [6] = 1'b0;
   assign \FB_filter[1][1] [5] = 1'b0;
   assign \FB_filter[1][1] [4] = 1'b0;
   assign \FB_filter[1][1] [3] = 1'b0;
   assign \FB_filter[1][1] [2] = 1'b0;
   assign \FB_filter[1][1] [1] = 1'b0;
   assign \FB_filter[1][1] [0] = 1'b0;
   assign \FB_filter[1][2] [15] = 1'b0;
   assign \FB_filter[1][2] [14] = 1'b0;
   assign \FB_filter[1][2] [13] = 1'b0;
   assign \FB_filter[1][2] [12] = 1'b0;
   assign \FB_filter[1][2] [11] = 1'b0;
   assign \FB_filter[1][2] [10] = 1'b0;
   assign \FB_filter[1][2] [9] = 1'b0;
   assign \FB_filter[1][2] [8] = 1'b0;
   assign \FB_filter[1][2] [7] = 1'b0;
   assign \FB_filter[1][2] [6] = 1'b0;
   assign \FB_filter[1][2] [5] = 1'b0;
   assign \FB_filter[1][2] [4] = 1'b0;
   assign \FB_filter[1][2] [3] = 1'b0;
   assign \FB_filter[1][2] [2] = 1'b0;
   assign \FB_filter[1][2] [1] = 1'b0;
   assign \FB_filter[1][2] [0] = 1'b0;
   assign \FB_filter[1][3] [15] = 1'b0;
   assign \FB_filter[1][3] [14] = 1'b0;
   assign \FB_filter[1][3] [13] = 1'b0;
   assign \FB_filter[1][3] [12] = 1'b0;
   assign \FB_filter[1][3] [11] = 1'b0;
   assign \FB_filter[1][3] [10] = 1'b0;
   assign \FB_filter[1][3] [9] = 1'b0;
   assign \FB_filter[1][3] [8] = 1'b0;
   assign \FB_filter[1][3] [7] = 1'b0;
   assign \FB_filter[1][3] [6] = 1'b0;
   assign \FB_filter[1][3] [5] = 1'b0;
   assign \FB_filter[1][3] [4] = 1'b0;
   assign \FB_filter[1][3] [3] = 1'b0;
   assign \FB_filter[1][3] [2] = 1'b0;
   assign \FB_filter[1][3] [1] = 1'b0;
   assign \FB_filter[1][3] [0] = 1'b0;
   assign \FB_filter[1][4] [15] = 1'b0;
   assign \FB_filter[1][4] [14] = 1'b0;
   assign \FB_filter[1][4] [13] = 1'b0;
   assign \FB_filter[1][4] [12] = 1'b0;
   assign \FB_filter[1][4] [11] = 1'b0;
   assign \FB_filter[1][4] [10] = 1'b0;
   assign \FB_filter[1][4] [9] = 1'b0;
   assign \FB_filter[1][4] [8] = 1'b0;
   assign \FB_filter[1][4] [7] = 1'b0;
   assign \FB_filter[1][4] [6] = 1'b0;
   assign \FB_filter[1][4] [5] = 1'b0;
   assign \FB_filter[1][4] [4] = 1'b0;
   assign \FB_filter[1][4] [3] = 1'b0;
   assign \FB_filter[1][4] [2] = 1'b0;
   assign \FB_filter[1][4] [1] = 1'b0;
   assign \FB_filter[1][4] [0] = 1'b0;
   assign \FB_filter[2][0] [15] = 1'b0;
   assign \FB_filter[2][0] [14] = 1'b0;
   assign \FB_filter[2][0] [13] = 1'b0;
   assign \FB_filter[2][0] [12] = 1'b0;
   assign \FB_filter[2][0] [11] = 1'b0;
   assign \FB_filter[2][0] [10] = 1'b0;
   assign \FB_filter[2][0] [9] = 1'b0;
   assign \FB_filter[2][0] [8] = 1'b0;
   assign \FB_filter[2][0] [7] = 1'b0;
   assign \FB_filter[2][0] [6] = 1'b0;
   assign \FB_filter[2][0] [5] = 1'b0;
   assign \FB_filter[2][0] [4] = 1'b0;
   assign \FB_filter[2][0] [3] = 1'b0;
   assign \FB_filter[2][0] [2] = 1'b0;
   assign \FB_filter[2][0] [1] = 1'b0;
   assign \FB_filter[2][0] [0] = 1'b0;
   assign \FB_filter[2][1] [15] = 1'b0;
   assign \FB_filter[2][1] [14] = 1'b0;
   assign \FB_filter[2][1] [13] = 1'b0;
   assign \FB_filter[2][1] [12] = 1'b0;
   assign \FB_filter[2][1] [11] = 1'b0;
   assign \FB_filter[2][1] [10] = 1'b0;
   assign \FB_filter[2][1] [9] = 1'b0;
   assign \FB_filter[2][1] [8] = 1'b0;
   assign \FB_filter[2][1] [7] = 1'b0;
   assign \FB_filter[2][1] [6] = 1'b0;
   assign \FB_filter[2][1] [5] = 1'b0;
   assign \FB_filter[2][1] [4] = 1'b0;
   assign \FB_filter[2][1] [3] = 1'b0;
   assign \FB_filter[2][1] [2] = 1'b0;
   assign \FB_filter[2][1] [1] = 1'b0;
   assign \FB_filter[2][1] [0] = 1'b0;
   assign \FB_filter[2][2] [15] = 1'b0;
   assign \FB_filter[2][2] [14] = 1'b0;
   assign \FB_filter[2][2] [13] = 1'b0;
   assign \FB_filter[2][2] [12] = 1'b0;
   assign \FB_filter[2][2] [11] = 1'b0;
   assign \FB_filter[2][2] [10] = 1'b0;
   assign \FB_filter[2][2] [9] = 1'b0;
   assign \FB_filter[2][2] [8] = 1'b0;
   assign \FB_filter[2][2] [7] = 1'b0;
   assign \FB_filter[2][2] [6] = 1'b0;
   assign \FB_filter[2][2] [5] = 1'b0;
   assign \FB_filter[2][2] [4] = 1'b0;
   assign \FB_filter[2][2] [3] = 1'b0;
   assign \FB_filter[2][2] [2] = 1'b0;
   assign \FB_filter[2][2] [1] = 1'b0;
   assign \FB_filter[2][2] [0] = 1'b0;
   assign \FB_filter[2][3] [15] = 1'b0;
   assign \FB_filter[2][3] [14] = 1'b0;
   assign \FB_filter[2][3] [13] = 1'b0;
   assign \FB_filter[2][3] [12] = 1'b0;
   assign \FB_filter[2][3] [11] = 1'b0;
   assign \FB_filter[2][3] [10] = 1'b0;
   assign \FB_filter[2][3] [9] = 1'b0;
   assign \FB_filter[2][3] [8] = 1'b0;
   assign \FB_filter[2][3] [7] = 1'b0;
   assign \FB_filter[2][3] [6] = 1'b0;
   assign \FB_filter[2][3] [5] = 1'b0;
   assign \FB_filter[2][3] [4] = 1'b0;
   assign \FB_filter[2][3] [3] = 1'b0;
   assign \FB_filter[2][3] [2] = 1'b0;
   assign \FB_filter[2][3] [1] = 1'b0;
   assign \FB_filter[2][3] [0] = 1'b0;
   assign \FB_filter[2][4] [15] = 1'b0;
   assign \FB_filter[2][4] [14] = 1'b0;
   assign \FB_filter[2][4] [13] = 1'b0;
   assign \FB_filter[2][4] [12] = 1'b0;
   assign \FB_filter[2][4] [11] = 1'b0;
   assign \FB_filter[2][4] [10] = 1'b0;
   assign \FB_filter[2][4] [9] = 1'b0;
   assign \FB_filter[2][4] [8] = 1'b0;
   assign \FB_filter[2][4] [7] = 1'b0;
   assign \FB_filter[2][4] [6] = 1'b0;
   assign \FB_filter[2][4] [5] = 1'b0;
   assign \FB_filter[2][4] [4] = 1'b0;
   assign \FB_filter[2][4] [3] = 1'b0;
   assign \FB_filter[2][4] [2] = 1'b0;
   assign \FB_filter[2][4] [1] = 1'b0;
   assign \FB_filter[2][4] [0] = 1'b0;
   assign \FB_filter[3][0] [15] = 1'b0;
   assign \FB_filter[3][0] [14] = 1'b0;
   assign \FB_filter[3][0] [13] = 1'b0;
   assign \FB_filter[3][0] [12] = 1'b0;
   assign \FB_filter[3][0] [11] = 1'b0;
   assign \FB_filter[3][0] [10] = 1'b0;
   assign \FB_filter[3][0] [9] = 1'b0;
   assign \FB_filter[3][0] [8] = 1'b0;
   assign \FB_filter[3][0] [7] = 1'b0;
   assign \FB_filter[3][0] [6] = 1'b0;
   assign \FB_filter[3][0] [5] = 1'b0;
   assign \FB_filter[3][0] [4] = 1'b0;
   assign \FB_filter[3][0] [3] = 1'b0;
   assign \FB_filter[3][0] [2] = 1'b0;
   assign \FB_filter[3][0] [1] = 1'b0;
   assign \FB_filter[3][0] [0] = 1'b0;
   assign \FB_filter[3][1] [15] = 1'b0;
   assign \FB_filter[3][1] [14] = 1'b0;
   assign \FB_filter[3][1] [13] = 1'b0;
   assign \FB_filter[3][1] [12] = 1'b0;
   assign \FB_filter[3][1] [11] = 1'b0;
   assign \FB_filter[3][1] [10] = 1'b0;
   assign \FB_filter[3][1] [9] = 1'b0;
   assign \FB_filter[3][1] [8] = 1'b0;
   assign \FB_filter[3][1] [7] = 1'b0;
   assign \FB_filter[3][1] [6] = 1'b0;
   assign \FB_filter[3][1] [5] = 1'b0;
   assign \FB_filter[3][1] [4] = 1'b0;
   assign \FB_filter[3][1] [3] = 1'b0;
   assign \FB_filter[3][1] [2] = 1'b0;
   assign \FB_filter[3][1] [1] = 1'b0;
   assign \FB_filter[3][1] [0] = 1'b0;
   assign \FB_filter[3][2] [15] = 1'b0;
   assign \FB_filter[3][2] [14] = 1'b0;
   assign \FB_filter[3][2] [13] = 1'b0;
   assign \FB_filter[3][2] [12] = 1'b0;
   assign \FB_filter[3][2] [11] = 1'b0;
   assign \FB_filter[3][2] [10] = 1'b0;
   assign \FB_filter[3][2] [9] = 1'b0;
   assign \FB_filter[3][2] [8] = 1'b0;
   assign \FB_filter[3][2] [7] = 1'b0;
   assign \FB_filter[3][2] [6] = 1'b0;
   assign \FB_filter[3][2] [5] = 1'b0;
   assign \FB_filter[3][2] [4] = 1'b0;
   assign \FB_filter[3][2] [3] = 1'b0;
   assign \FB_filter[3][2] [2] = 1'b0;
   assign \FB_filter[3][2] [1] = 1'b0;
   assign \FB_filter[3][2] [0] = 1'b0;
   assign \FB_filter[3][3] [15] = 1'b0;
   assign \FB_filter[3][3] [14] = 1'b0;
   assign \FB_filter[3][3] [13] = 1'b0;
   assign \FB_filter[3][3] [12] = 1'b0;
   assign \FB_filter[3][3] [11] = 1'b0;
   assign \FB_filter[3][3] [10] = 1'b0;
   assign \FB_filter[3][3] [9] = 1'b0;
   assign \FB_filter[3][3] [8] = 1'b0;
   assign \FB_filter[3][3] [7] = 1'b0;
   assign \FB_filter[3][3] [6] = 1'b0;
   assign \FB_filter[3][3] [5] = 1'b0;
   assign \FB_filter[3][3] [4] = 1'b0;
   assign \FB_filter[3][3] [3] = 1'b0;
   assign \FB_filter[3][3] [2] = 1'b0;
   assign \FB_filter[3][3] [1] = 1'b0;
   assign \FB_filter[3][3] [0] = 1'b0;
   assign \FB_filter[3][4] [15] = 1'b0;
   assign \FB_filter[3][4] [14] = 1'b0;
   assign \FB_filter[3][4] [13] = 1'b0;
   assign \FB_filter[3][4] [12] = 1'b0;
   assign \FB_filter[3][4] [11] = 1'b0;
   assign \FB_filter[3][4] [10] = 1'b0;
   assign \FB_filter[3][4] [9] = 1'b0;
   assign \FB_filter[3][4] [8] = 1'b0;
   assign \FB_filter[3][4] [7] = 1'b0;
   assign \FB_filter[3][4] [6] = 1'b0;
   assign \FB_filter[3][4] [5] = 1'b0;
   assign \FB_filter[3][4] [4] = 1'b0;
   assign \FB_filter[3][4] [3] = 1'b0;
   assign \FB_filter[3][4] [2] = 1'b0;
   assign \FB_filter[3][4] [1] = 1'b0;
   assign \FB_filter[3][4] [0] = 1'b0;
   assign \FB_filter[4][0] [15] = 1'b0;
   assign \FB_filter[4][0] [14] = 1'b0;
   assign \FB_filter[4][0] [13] = 1'b0;
   assign \FB_filter[4][0] [12] = 1'b0;
   assign \FB_filter[4][0] [11] = 1'b0;
   assign \FB_filter[4][0] [10] = 1'b0;
   assign \FB_filter[4][0] [9] = 1'b0;
   assign \FB_filter[4][0] [8] = 1'b0;
   assign \FB_filter[4][0] [7] = 1'b0;
   assign \FB_filter[4][0] [6] = 1'b0;
   assign \FB_filter[4][0] [5] = 1'b0;
   assign \FB_filter[4][0] [4] = 1'b0;
   assign \FB_filter[4][0] [3] = 1'b0;
   assign \FB_filter[4][0] [2] = 1'b0;
   assign \FB_filter[4][0] [1] = 1'b0;
   assign \FB_filter[4][0] [0] = 1'b0;
   assign \FB_filter[4][1] [15] = 1'b0;
   assign \FB_filter[4][1] [14] = 1'b0;
   assign \FB_filter[4][1] [13] = 1'b0;
   assign \FB_filter[4][1] [12] = 1'b0;
   assign \FB_filter[4][1] [11] = 1'b0;
   assign \FB_filter[4][1] [10] = 1'b0;
   assign \FB_filter[4][1] [9] = 1'b0;
   assign \FB_filter[4][1] [8] = 1'b0;
   assign \FB_filter[4][1] [7] = 1'b0;
   assign \FB_filter[4][1] [6] = 1'b0;
   assign \FB_filter[4][1] [5] = 1'b0;
   assign \FB_filter[4][1] [4] = 1'b0;
   assign \FB_filter[4][1] [3] = 1'b0;
   assign \FB_filter[4][1] [2] = 1'b0;
   assign \FB_filter[4][1] [1] = 1'b0;
   assign \FB_filter[4][1] [0] = 1'b0;
   assign \FB_filter[4][2] [15] = 1'b0;
   assign \FB_filter[4][2] [14] = 1'b0;
   assign \FB_filter[4][2] [13] = 1'b0;
   assign \FB_filter[4][2] [12] = 1'b0;
   assign \FB_filter[4][2] [11] = 1'b0;
   assign \FB_filter[4][2] [10] = 1'b0;
   assign \FB_filter[4][2] [9] = 1'b0;
   assign \FB_filter[4][2] [8] = 1'b0;
   assign \FB_filter[4][2] [7] = 1'b0;
   assign \FB_filter[4][2] [6] = 1'b0;
   assign \FB_filter[4][2] [5] = 1'b0;
   assign \FB_filter[4][2] [4] = 1'b0;
   assign \FB_filter[4][2] [3] = 1'b0;
   assign \FB_filter[4][2] [2] = 1'b0;
   assign \FB_filter[4][2] [1] = 1'b0;
   assign \FB_filter[4][2] [0] = 1'b0;
   assign \FB_filter[4][3] [15] = 1'b0;
   assign \FB_filter[4][3] [14] = 1'b0;
   assign \FB_filter[4][3] [13] = 1'b0;
   assign \FB_filter[4][3] [12] = 1'b0;
   assign \FB_filter[4][3] [11] = 1'b0;
   assign \FB_filter[4][3] [10] = 1'b0;
   assign \FB_filter[4][3] [9] = 1'b0;
   assign \FB_filter[4][3] [8] = 1'b0;
   assign \FB_filter[4][3] [7] = 1'b0;
   assign \FB_filter[4][3] [6] = 1'b0;
   assign \FB_filter[4][3] [5] = 1'b0;
   assign \FB_filter[4][3] [4] = 1'b0;
   assign \FB_filter[4][3] [3] = 1'b0;
   assign \FB_filter[4][3] [2] = 1'b0;
   assign \FB_filter[4][3] [1] = 1'b0;
   assign \FB_filter[4][3] [0] = 1'b0;
   assign \FB_filter[4][4] [15] = 1'b0;
   assign \FB_filter[4][4] [14] = 1'b0;
   assign \FB_filter[4][4] [13] = 1'b0;
   assign \FB_filter[4][4] [12] = 1'b0;
   assign \FB_filter[4][4] [11] = 1'b0;
   assign \FB_filter[4][4] [10] = 1'b0;
   assign \FB_filter[4][4] [9] = 1'b0;
   assign \FB_filter[4][4] [8] = 1'b0;
   assign \FB_filter[4][4] [7] = 1'b0;
   assign \FB_filter[4][4] [6] = 1'b0;
   assign \FB_filter[4][4] [5] = 1'b0;
   assign \FB_filter[4][4] [4] = 1'b0;
   assign \FB_filter[4][4] [3] = 1'b0;
   assign \FB_filter[4][4] [2] = 1'b0;
   assign \FB_filter[4][4] [1] = 1'b0;
   assign \FB_filter[4][4] [0] = 1'b0;
   assign FB_index_filter[15] = 1'b0;
   assign FB_index_filter[14] = 1'b0;
   assign FB_index_filter[13] = 1'b0;
   assign FB_index_filter[12] = 1'b0;
   assign FB_index_filter[11] = 1'b0;
   assign FB_index_filter[10] = 1'b0;
   assign FB_index_filter[9] = 1'b0;
   assign FB_index_filter[8] = 1'b0;
   assign FB_index_filter[7] = 1'b0;
   assign FB_index_filter[6] = 1'b0;
   assign FB_index_filter[5] = 1'b0;
   assign FB_index_filter[4] = 1'b0;
   assign FB_index_filter[3] = 1'b0;
   assign FB_index_filter[2] = 1'b0;
   assign FB_index_filter[1] = 1'b0;
   assign FB_index_filter[0] = 1'b0;

   datapath__0_73 i_1_14 (.p_0({1'b0, uc_0, uc_1, 1'b0, 1'b0, RAM_finish}), 
      .p_1({n_1_52, n_1_51, n_1_50, n_1_49, n_1_48, n_1_47, n_1_46, n_1_45, 
      n_1_28, n_1_27, n_1_26, n_1_25, n_1_24, n_1_23, n_1_22, n_1_21}), 
      .inner_address({n_1_44, n_1_43, n_1_42, n_1_41, n_1_40, n_1_39, n_1_38, 
      n_1_37, n_1_36, n_1_35, n_1_34, n_1_33, n_1_32, n_1_31, n_1_30, n_1_29}));
   HA_X1 i_1_0_0 (.A(biasCounter[2]), .B(n_1_0_3), .CO(n_1_0_1), .S());
   HA_X1 i_1_0_1 (.A(biasCounter[1]), .B(biasCounter[0]), .CO(n_1_0_0), .S(
      n_1_0_4));
   HA_X1 i_1_0_2 (.A(biasCounter[2]), .B(n_1_0_0), .CO(n_1_0_2), .S(n_1_0_5));
   NOR2_X1 i_1_0_3 (.A1(biasCounter[0]), .A2(n_1_0_44), .ZN(n_1_0));
   AND2_X1 i_1_0_4 (.A1(n_1_0_43), .A2(n_1_0_4), .ZN(n_1_1));
   AND2_X1 i_1_0_5 (.A1(n_1_0_43), .A2(n_1_0_5), .ZN(n_1_2));
   OAI21_X1 i_1_0_6 (.A(n_1_0_6), .B1(n_1_0_2), .B2(n_1_0_54), .ZN(n_1_3));
   NAND3_X1 i_1_0_7 (.A1(n_1_0_54), .A2(n_1_0_50), .A3(n_1_0_2), .ZN(n_1_0_6));
   AOI21_X1 i_1_0_8 (.A(n_1_0_47), .B1(n_1_0_43), .B2(n_1_0_53), .ZN(n_1_4));
   NOR2_X1 i_1_0_9 (.A1(n_1_0_53), .A2(n_1_0_45), .ZN(n_1_5));
   INV_X1 i_1_0_10 (.A(n_1_0_7), .ZN(n_1_77));
   AOI22_X1 i_1_0_11 (.A1(n_1_0_24), .A2(address[0]), .B1(inner_address[0]), 
      .B2(n_1_0_23), .ZN(n_1_0_7));
   INV_X1 i_1_0_12 (.A(n_1_0_8), .ZN(n_1_6));
   AOI22_X1 i_1_0_13 (.A1(n_1_0_24), .A2(address[1]), .B1(inner_address[1]), 
      .B2(n_1_0_23), .ZN(n_1_0_8));
   INV_X1 i_1_0_14 (.A(n_1_0_9), .ZN(n_1_7));
   AOI22_X1 i_1_0_15 (.A1(n_1_0_24), .A2(address[2]), .B1(inner_address[2]), 
      .B2(n_1_0_23), .ZN(n_1_0_9));
   INV_X1 i_1_0_16 (.A(n_1_0_10), .ZN(n_1_8));
   AOI22_X1 i_1_0_17 (.A1(n_1_0_24), .A2(address[3]), .B1(inner_address[3]), 
      .B2(n_1_0_23), .ZN(n_1_0_10));
   INV_X1 i_1_0_18 (.A(n_1_0_11), .ZN(n_1_9));
   AOI22_X1 i_1_0_19 (.A1(n_1_0_24), .A2(address[4]), .B1(inner_address[4]), 
      .B2(n_1_0_23), .ZN(n_1_0_11));
   INV_X1 i_1_0_20 (.A(n_1_0_12), .ZN(n_1_10));
   AOI22_X1 i_1_0_21 (.A1(n_1_0_24), .A2(address[5]), .B1(inner_address[5]), 
      .B2(n_1_0_23), .ZN(n_1_0_12));
   INV_X1 i_1_0_22 (.A(n_1_0_13), .ZN(n_1_11));
   AOI22_X1 i_1_0_23 (.A1(n_1_0_24), .A2(address[6]), .B1(inner_address[6]), 
      .B2(n_1_0_23), .ZN(n_1_0_13));
   INV_X1 i_1_0_24 (.A(n_1_0_14), .ZN(n_1_12));
   AOI22_X1 i_1_0_25 (.A1(n_1_0_24), .A2(address[7]), .B1(inner_address[7]), 
      .B2(n_1_0_23), .ZN(n_1_0_14));
   INV_X1 i_1_0_26 (.A(n_1_0_15), .ZN(n_1_13));
   AOI22_X1 i_1_0_27 (.A1(n_1_0_24), .A2(address[8]), .B1(inner_address[8]), 
      .B2(n_1_0_23), .ZN(n_1_0_15));
   INV_X1 i_1_0_28 (.A(n_1_0_16), .ZN(n_1_14));
   AOI22_X1 i_1_0_29 (.A1(n_1_0_24), .A2(address[9]), .B1(inner_address[9]), 
      .B2(n_1_0_23), .ZN(n_1_0_16));
   INV_X1 i_1_0_30 (.A(n_1_0_17), .ZN(n_1_15));
   AOI22_X1 i_1_0_31 (.A1(n_1_0_24), .A2(address[10]), .B1(inner_address[10]), 
      .B2(n_1_0_23), .ZN(n_1_0_17));
   INV_X1 i_1_0_32 (.A(n_1_0_18), .ZN(n_1_16));
   AOI22_X1 i_1_0_33 (.A1(n_1_0_24), .A2(address[11]), .B1(inner_address[11]), 
      .B2(n_1_0_23), .ZN(n_1_0_18));
   INV_X1 i_1_0_34 (.A(n_1_0_19), .ZN(n_1_17));
   AOI22_X1 i_1_0_35 (.A1(n_1_0_24), .A2(address[12]), .B1(inner_address[12]), 
      .B2(n_1_0_23), .ZN(n_1_0_19));
   INV_X1 i_1_0_36 (.A(n_1_0_20), .ZN(n_1_18));
   AOI22_X1 i_1_0_37 (.A1(n_1_0_24), .A2(address[13]), .B1(inner_address[13]), 
      .B2(n_1_0_23), .ZN(n_1_0_20));
   INV_X1 i_1_0_38 (.A(n_1_0_21), .ZN(n_1_19));
   AOI22_X1 i_1_0_39 (.A1(n_1_0_24), .A2(address[14]), .B1(inner_address[14]), 
      .B2(n_1_0_23), .ZN(n_1_0_21));
   INV_X1 i_1_0_40 (.A(n_1_0_22), .ZN(n_1_20));
   AOI22_X1 i_1_0_41 (.A1(n_1_0_24), .A2(address[15]), .B1(inner_address[15]), 
      .B2(n_1_0_23), .ZN(n_1_0_22));
   AOI21_X1 i_1_0_42 (.A(n_1_0_52), .B1(read_write_filter_bias[0]), .B2(n_1_0_42), 
      .ZN(n_1_0_23));
   OAI21_X1 i_1_0_43 (.A(n_1_0_25), .B1(read_write_filter_bias[0]), .B2(
      read_write_filter_bias[1]), .ZN(n_1_0_24));
   NAND2_X1 i_1_0_44 (.A1(n_1_0_48), .A2(n_1_0_42), .ZN(n_1_0_25));
   INV_X1 i_1_0_45 (.A(n_1_0_26), .ZN(n_1_61));
   AOI22_X1 i_1_0_46 (.A1(inner_address[0]), .A2(n_1_0_49), .B1(n_1_0_48), 
      .B2(n_1_29), .ZN(n_1_0_26));
   INV_X1 i_1_0_47 (.A(n_1_0_27), .ZN(n_1_62));
   AOI22_X1 i_1_0_48 (.A1(inner_address[1]), .A2(n_1_0_49), .B1(n_1_0_48), 
      .B2(n_1_30), .ZN(n_1_0_27));
   INV_X1 i_1_0_49 (.A(n_1_0_28), .ZN(n_1_63));
   AOI22_X1 i_1_0_50 (.A1(inner_address[2]), .A2(n_1_0_49), .B1(n_1_0_48), 
      .B2(n_1_31), .ZN(n_1_0_28));
   INV_X1 i_1_0_51 (.A(n_1_0_29), .ZN(n_1_64));
   AOI22_X1 i_1_0_52 (.A1(inner_address[3]), .A2(n_1_0_49), .B1(n_1_0_48), 
      .B2(n_1_32), .ZN(n_1_0_29));
   INV_X1 i_1_0_53 (.A(n_1_0_30), .ZN(n_1_65));
   AOI22_X1 i_1_0_54 (.A1(inner_address[4]), .A2(n_1_0_49), .B1(n_1_0_48), 
      .B2(n_1_33), .ZN(n_1_0_30));
   INV_X1 i_1_0_55 (.A(n_1_0_31), .ZN(n_1_66));
   AOI22_X1 i_1_0_56 (.A1(inner_address[5]), .A2(n_1_0_49), .B1(n_1_0_48), 
      .B2(n_1_34), .ZN(n_1_0_31));
   INV_X1 i_1_0_57 (.A(n_1_0_32), .ZN(n_1_67));
   AOI22_X1 i_1_0_58 (.A1(inner_address[6]), .A2(n_1_0_49), .B1(n_1_0_48), 
      .B2(n_1_35), .ZN(n_1_0_32));
   INV_X1 i_1_0_59 (.A(n_1_0_33), .ZN(n_1_68));
   AOI22_X1 i_1_0_60 (.A1(inner_address[7]), .A2(n_1_0_49), .B1(n_1_0_48), 
      .B2(n_1_36), .ZN(n_1_0_33));
   INV_X1 i_1_0_61 (.A(n_1_0_34), .ZN(n_1_69));
   AOI22_X1 i_1_0_62 (.A1(inner_address[8]), .A2(n_1_0_49), .B1(n_1_0_48), 
      .B2(n_1_37), .ZN(n_1_0_34));
   INV_X1 i_1_0_63 (.A(n_1_0_35), .ZN(n_1_70));
   AOI22_X1 i_1_0_64 (.A1(inner_address[9]), .A2(n_1_0_49), .B1(n_1_0_48), 
      .B2(n_1_38), .ZN(n_1_0_35));
   INV_X1 i_1_0_65 (.A(n_1_0_36), .ZN(n_1_71));
   AOI22_X1 i_1_0_66 (.A1(inner_address[10]), .A2(n_1_0_49), .B1(n_1_0_48), 
      .B2(n_1_39), .ZN(n_1_0_36));
   INV_X1 i_1_0_67 (.A(n_1_0_37), .ZN(n_1_72));
   AOI22_X1 i_1_0_68 (.A1(inner_address[11]), .A2(n_1_0_49), .B1(n_1_0_48), 
      .B2(n_1_40), .ZN(n_1_0_37));
   INV_X1 i_1_0_69 (.A(n_1_0_38), .ZN(n_1_73));
   AOI22_X1 i_1_0_70 (.A1(inner_address[12]), .A2(n_1_0_49), .B1(n_1_0_48), 
      .B2(n_1_41), .ZN(n_1_0_38));
   INV_X1 i_1_0_71 (.A(n_1_0_39), .ZN(n_1_74));
   AOI22_X1 i_1_0_72 (.A1(inner_address[13]), .A2(n_1_0_49), .B1(n_1_0_48), 
      .B2(n_1_42), .ZN(n_1_0_39));
   INV_X1 i_1_0_73 (.A(n_1_0_40), .ZN(n_1_75));
   AOI22_X1 i_1_0_74 (.A1(inner_address[14]), .A2(n_1_0_49), .B1(n_1_0_48), 
      .B2(n_1_43), .ZN(n_1_0_40));
   INV_X1 i_1_0_75 (.A(n_1_0_41), .ZN(n_1_76));
   AOI22_X1 i_1_0_76 (.A1(inner_address[15]), .A2(n_1_0_49), .B1(n_1_0_48), 
      .B2(n_1_44), .ZN(n_1_0_41));
   MUX2_X1 i_1_0_77 (.A(inner_address[0]), .B(address[0]), .S(n_1_0_42), 
      .Z(n_1_21));
   MUX2_X1 i_1_0_78 (.A(inner_address[1]), .B(address[1]), .S(n_1_0_42), 
      .Z(n_1_22));
   MUX2_X1 i_1_0_79 (.A(inner_address[2]), .B(address[2]), .S(n_1_0_42), 
      .Z(n_1_23));
   MUX2_X1 i_1_0_80 (.A(inner_address[3]), .B(address[3]), .S(n_1_0_42), 
      .Z(n_1_24));
   MUX2_X1 i_1_0_81 (.A(inner_address[4]), .B(address[4]), .S(n_1_0_42), 
      .Z(n_1_25));
   MUX2_X1 i_1_0_82 (.A(inner_address[5]), .B(address[5]), .S(n_1_0_42), 
      .Z(n_1_26));
   MUX2_X1 i_1_0_83 (.A(inner_address[6]), .B(address[6]), .S(n_1_0_42), 
      .Z(n_1_27));
   MUX2_X1 i_1_0_84 (.A(inner_address[7]), .B(address[7]), .S(n_1_0_42), 
      .Z(n_1_28));
   MUX2_X1 i_1_0_85 (.A(inner_address[8]), .B(address[8]), .S(n_1_0_42), 
      .Z(n_1_45));
   MUX2_X1 i_1_0_86 (.A(inner_address[9]), .B(address[9]), .S(n_1_0_42), 
      .Z(n_1_46));
   MUX2_X1 i_1_0_87 (.A(inner_address[10]), .B(address[10]), .S(n_1_0_42), 
      .Z(n_1_47));
   MUX2_X1 i_1_0_88 (.A(inner_address[11]), .B(address[11]), .S(n_1_0_42), 
      .Z(n_1_48));
   MUX2_X1 i_1_0_89 (.A(inner_address[12]), .B(address[12]), .S(n_1_0_42), 
      .Z(n_1_49));
   MUX2_X1 i_1_0_90 (.A(inner_address[13]), .B(address[13]), .S(n_1_0_42), 
      .Z(n_1_50));
   MUX2_X1 i_1_0_91 (.A(inner_address[14]), .B(address[14]), .S(n_1_0_42), 
      .Z(n_1_51));
   MUX2_X1 i_1_0_92 (.A(inner_address[15]), .B(address[15]), .S(n_1_0_42), 
      .Z(n_1_52));
   NOR3_X1 i_1_0_93 (.A1(n_1_0_3), .A2(biasCounter[2]), .A3(biasCounter[31]), 
      .ZN(n_1_0_42));
   OR2_X1 i_1_0_94 (.A1(biasCounter[1]), .A2(biasCounter[0]), .ZN(n_1_0_3));
   OAI21_X1 i_1_0_95 (.A(n_1_0_45), .B1(n_1_0_47), .B2(n_1_0_44), .ZN(n_1_54));
   NOR2_X1 i_1_0_96 (.A1(n_1_0_47), .A2(n_1_0_44), .ZN(n_1_53));
   NAND2_X1 i_1_0_97 (.A1(n_1_0_54), .A2(n_1_0_1), .ZN(n_1_0_43));
   NOR2_X1 i_1_0_98 (.A1(n_1_0_50), .A2(biasCounter[31]), .ZN(n_1_0_44));
   NAND3_X1 i_1_0_99 (.A1(n_1_0_52), .A2(n_1_0_51), .A3(start), .ZN(n_1_0_45));
   NOR2_X1 i_1_0_100 (.A1(n_1_0_47), .A2(n_1_0_46), .ZN(n_1_78));
   NAND4_X1 i_1_0_101 (.A1(n_1_0_54), .A2(n_1_0_50), .A3(RAM_finish), .A4(
      biasCounter[2]), .ZN(n_1_0_46));
   NAND2_X1 i_1_0_102 (.A1(start), .A2(n_1_0_48), .ZN(n_1_0_47));
   NOR2_X1 i_1_0_103 (.A1(n_1_0_52), .A2(n_1_0_51), .ZN(n_1_0_48));
   NOR3_X1 i_1_0_104 (.A1(n_1_0_53), .A2(n_1_0_52), .A3(
      read_write_filter_bias[0]), .ZN(n_1_55));
   NOR2_X1 i_1_0_105 (.A1(n_1_0_52), .A2(read_write_filter_bias[0]), .ZN(
      n_1_0_49));
   INV_X1 i_1_0_106 (.A(n_1_0_1), .ZN(n_1_0_50));
   INV_X1 i_1_0_107 (.A(read_write_filter_bias[0]), .ZN(n_1_0_51));
   INV_X1 i_1_0_108 (.A(read_write_filter_bias[1]), .ZN(n_1_0_52));
   INV_X1 i_1_0_109 (.A(RAM_finish), .ZN(n_1_0_53));
   INV_X1 i_1_0_110 (.A(biasCounter[31]), .ZN(n_1_0_54));
   DFF_X1 \CNN_output_data_reg[4][4][15]  (.D(\RAM_input_data[4][4] [15]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][4] [15]), .QN());
   DFF_X1 \CNN_output_data_reg[4][4][14]  (.D(\RAM_input_data[4][4] [14]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][4] [14]), .QN());
   DFF_X1 \CNN_output_data_reg[4][4][13]  (.D(\RAM_input_data[4][4] [13]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][4] [13]), .QN());
   DFF_X1 \CNN_output_data_reg[4][4][12]  (.D(\RAM_input_data[4][4] [12]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][4] [12]), .QN());
   DFF_X1 \CNN_output_data_reg[4][4][11]  (.D(\RAM_input_data[4][4] [11]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][4] [11]), .QN());
   DFF_X1 \CNN_output_data_reg[4][4][10]  (.D(\RAM_input_data[4][4] [10]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][4] [10]), .QN());
   DFF_X1 \CNN_output_data_reg[4][4][9]  (.D(\RAM_input_data[4][4] [9]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][4] [9]), .QN());
   DFF_X1 \CNN_output_data_reg[4][4][8]  (.D(\RAM_input_data[4][4] [8]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][4] [8]), .QN());
   DFF_X1 \CNN_output_data_reg[4][4][7]  (.D(\RAM_input_data[4][4] [7]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][4] [7]), .QN());
   DFF_X1 \CNN_output_data_reg[4][4][6]  (.D(\RAM_input_data[4][4] [6]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][4] [6]), .QN());
   DFF_X1 \CNN_output_data_reg[4][4][5]  (.D(\RAM_input_data[4][4] [5]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][4] [5]), .QN());
   DFF_X1 \CNN_output_data_reg[4][4][4]  (.D(\RAM_input_data[4][4] [4]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][4] [4]), .QN());
   DFF_X1 \CNN_output_data_reg[4][4][3]  (.D(\RAM_input_data[4][4] [3]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][4] [3]), .QN());
   DFF_X1 \CNN_output_data_reg[4][4][2]  (.D(\RAM_input_data[4][4] [2]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][4] [2]), .QN());
   DFF_X1 \CNN_output_data_reg[4][4][1]  (.D(\RAM_input_data[4][4] [1]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][4] [1]), .QN());
   DFF_X1 \CNN_output_data_reg[4][4][0]  (.D(\RAM_input_data[4][4] [0]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][4] [0]), .QN());
   DFF_X1 \CNN_output_data_reg[4][3][15]  (.D(\RAM_input_data[4][3] [15]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][3] [15]), .QN());
   DFF_X1 \CNN_output_data_reg[4][3][14]  (.D(\RAM_input_data[4][3] [14]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][3] [14]), .QN());
   DFF_X1 \CNN_output_data_reg[4][3][13]  (.D(\RAM_input_data[4][3] [13]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][3] [13]), .QN());
   DFF_X1 \CNN_output_data_reg[4][3][12]  (.D(\RAM_input_data[4][3] [12]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][3] [12]), .QN());
   DFF_X1 \CNN_output_data_reg[4][3][11]  (.D(\RAM_input_data[4][3] [11]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][3] [11]), .QN());
   DFF_X1 \CNN_output_data_reg[4][3][10]  (.D(\RAM_input_data[4][3] [10]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][3] [10]), .QN());
   DFF_X1 \CNN_output_data_reg[4][3][9]  (.D(\RAM_input_data[4][3] [9]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][3] [9]), .QN());
   DFF_X1 \CNN_output_data_reg[4][3][8]  (.D(\RAM_input_data[4][3] [8]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][3] [8]), .QN());
   DFF_X1 \CNN_output_data_reg[4][3][7]  (.D(\RAM_input_data[4][3] [7]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][3] [7]), .QN());
   DFF_X1 \CNN_output_data_reg[4][3][6]  (.D(\RAM_input_data[4][3] [6]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][3] [6]), .QN());
   DFF_X1 \CNN_output_data_reg[4][3][5]  (.D(\RAM_input_data[4][3] [5]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][3] [5]), .QN());
   DFF_X1 \CNN_output_data_reg[4][3][4]  (.D(\RAM_input_data[4][3] [4]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][3] [4]), .QN());
   DFF_X1 \CNN_output_data_reg[4][3][3]  (.D(\RAM_input_data[4][3] [3]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][3] [3]), .QN());
   DFF_X1 \CNN_output_data_reg[4][3][2]  (.D(\RAM_input_data[4][3] [2]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][3] [2]), .QN());
   DFF_X1 \CNN_output_data_reg[4][3][1]  (.D(\RAM_input_data[4][3] [1]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][3] [1]), .QN());
   DFF_X1 \CNN_output_data_reg[4][3][0]  (.D(\RAM_input_data[4][3] [0]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][3] [0]), .QN());
   DFF_X1 \CNN_output_data_reg[4][2][15]  (.D(\RAM_input_data[4][2] [15]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][2] [15]), .QN());
   DFF_X1 \CNN_output_data_reg[4][2][14]  (.D(\RAM_input_data[4][2] [14]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][2] [14]), .QN());
   DFF_X1 \CNN_output_data_reg[4][2][13]  (.D(\RAM_input_data[4][2] [13]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][2] [13]), .QN());
   DFF_X1 \CNN_output_data_reg[4][2][12]  (.D(\RAM_input_data[4][2] [12]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][2] [12]), .QN());
   DFF_X1 \CNN_output_data_reg[4][2][11]  (.D(\RAM_input_data[4][2] [11]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][2] [11]), .QN());
   DFF_X1 \CNN_output_data_reg[4][2][10]  (.D(\RAM_input_data[4][2] [10]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][2] [10]), .QN());
   DFF_X1 \CNN_output_data_reg[4][2][9]  (.D(\RAM_input_data[4][2] [9]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][2] [9]), .QN());
   DFF_X1 \CNN_output_data_reg[4][2][8]  (.D(\RAM_input_data[4][2] [8]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][2] [8]), .QN());
   DFF_X1 \CNN_output_data_reg[4][2][7]  (.D(\RAM_input_data[4][2] [7]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][2] [7]), .QN());
   DFF_X1 \CNN_output_data_reg[4][2][6]  (.D(\RAM_input_data[4][2] [6]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][2] [6]), .QN());
   DFF_X1 \CNN_output_data_reg[4][2][5]  (.D(\RAM_input_data[4][2] [5]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][2] [5]), .QN());
   DFF_X1 \CNN_output_data_reg[4][2][4]  (.D(\RAM_input_data[4][2] [4]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][2] [4]), .QN());
   DFF_X1 \CNN_output_data_reg[4][2][3]  (.D(\RAM_input_data[4][2] [3]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][2] [3]), .QN());
   DFF_X1 \CNN_output_data_reg[4][2][2]  (.D(\RAM_input_data[4][2] [2]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][2] [2]), .QN());
   DFF_X1 \CNN_output_data_reg[4][2][1]  (.D(\RAM_input_data[4][2] [1]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][2] [1]), .QN());
   DFF_X1 \CNN_output_data_reg[4][2][0]  (.D(\RAM_input_data[4][2] [0]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][2] [0]), .QN());
   DFF_X1 \CNN_output_data_reg[4][1][15]  (.D(\RAM_input_data[4][1] [15]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][1] [15]), .QN());
   DFF_X1 \CNN_output_data_reg[4][1][14]  (.D(\RAM_input_data[4][1] [14]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][1] [14]), .QN());
   DFF_X1 \CNN_output_data_reg[4][1][13]  (.D(\RAM_input_data[4][1] [13]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][1] [13]), .QN());
   DFF_X1 \CNN_output_data_reg[4][1][12]  (.D(\RAM_input_data[4][1] [12]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][1] [12]), .QN());
   DFF_X1 \CNN_output_data_reg[4][1][11]  (.D(\RAM_input_data[4][1] [11]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][1] [11]), .QN());
   DFF_X1 \CNN_output_data_reg[4][1][10]  (.D(\RAM_input_data[4][1] [10]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][1] [10]), .QN());
   DFF_X1 \CNN_output_data_reg[4][1][9]  (.D(\RAM_input_data[4][1] [9]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][1] [9]), .QN());
   DFF_X1 \CNN_output_data_reg[4][1][8]  (.D(\RAM_input_data[4][1] [8]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][1] [8]), .QN());
   DFF_X1 \CNN_output_data_reg[4][1][7]  (.D(\RAM_input_data[4][1] [7]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][1] [7]), .QN());
   DFF_X1 \CNN_output_data_reg[4][1][6]  (.D(\RAM_input_data[4][1] [6]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][1] [6]), .QN());
   DFF_X1 \CNN_output_data_reg[4][1][5]  (.D(\RAM_input_data[4][1] [5]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][1] [5]), .QN());
   DFF_X1 \CNN_output_data_reg[4][1][4]  (.D(\RAM_input_data[4][1] [4]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][1] [4]), .QN());
   DFF_X1 \CNN_output_data_reg[4][1][3]  (.D(\RAM_input_data[4][1] [3]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][1] [3]), .QN());
   DFF_X1 \CNN_output_data_reg[4][1][2]  (.D(\RAM_input_data[4][1] [2]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][1] [2]), .QN());
   DFF_X1 \CNN_output_data_reg[4][1][1]  (.D(\RAM_input_data[4][1] [1]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][1] [1]), .QN());
   DFF_X1 \CNN_output_data_reg[4][1][0]  (.D(\RAM_input_data[4][1] [0]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][1] [0]), .QN());
   DFF_X1 \CNN_output_data_reg[4][0][15]  (.D(\RAM_input_data[4][0] [15]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][0] [15]), .QN());
   DFF_X1 \CNN_output_data_reg[4][0][14]  (.D(\RAM_input_data[4][0] [14]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][0] [14]), .QN());
   DFF_X1 \CNN_output_data_reg[4][0][13]  (.D(\RAM_input_data[4][0] [13]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][0] [13]), .QN());
   DFF_X1 \CNN_output_data_reg[4][0][12]  (.D(\RAM_input_data[4][0] [12]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][0] [12]), .QN());
   DFF_X1 \CNN_output_data_reg[4][0][11]  (.D(\RAM_input_data[4][0] [11]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][0] [11]), .QN());
   DFF_X1 \CNN_output_data_reg[4][0][10]  (.D(\RAM_input_data[4][0] [10]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][0] [10]), .QN());
   DFF_X1 \CNN_output_data_reg[4][0][9]  (.D(\RAM_input_data[4][0] [9]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][0] [9]), .QN());
   DFF_X1 \CNN_output_data_reg[4][0][8]  (.D(\RAM_input_data[4][0] [8]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][0] [8]), .QN());
   DFF_X1 \CNN_output_data_reg[4][0][7]  (.D(\RAM_input_data[4][0] [7]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][0] [7]), .QN());
   DFF_X1 \CNN_output_data_reg[4][0][6]  (.D(\RAM_input_data[4][0] [6]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][0] [6]), .QN());
   DFF_X1 \CNN_output_data_reg[4][0][5]  (.D(\RAM_input_data[4][0] [5]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][0] [5]), .QN());
   DFF_X1 \CNN_output_data_reg[4][0][4]  (.D(\RAM_input_data[4][0] [4]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][0] [4]), .QN());
   DFF_X1 \CNN_output_data_reg[4][0][3]  (.D(\RAM_input_data[4][0] [3]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][0] [3]), .QN());
   DFF_X1 \CNN_output_data_reg[4][0][2]  (.D(\RAM_input_data[4][0] [2]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][0] [2]), .QN());
   DFF_X1 \CNN_output_data_reg[4][0][1]  (.D(\RAM_input_data[4][0] [1]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][0] [1]), .QN());
   DFF_X1 \CNN_output_data_reg[4][0][0]  (.D(\RAM_input_data[4][0] [0]), 
      .CK(n_1_56), .Q(\CNN_output_data[4][0] [0]), .QN());
   DFF_X1 \CNN_output_data_reg[3][4][15]  (.D(\RAM_input_data[3][4] [15]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][4] [15]), .QN());
   DFF_X1 \CNN_output_data_reg[3][4][14]  (.D(\RAM_input_data[3][4] [14]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][4] [14]), .QN());
   DFF_X1 \CNN_output_data_reg[3][4][13]  (.D(\RAM_input_data[3][4] [13]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][4] [13]), .QN());
   DFF_X1 \CNN_output_data_reg[3][4][12]  (.D(\RAM_input_data[3][4] [12]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][4] [12]), .QN());
   DFF_X1 \CNN_output_data_reg[3][4][11]  (.D(\RAM_input_data[3][4] [11]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][4] [11]), .QN());
   DFF_X1 \CNN_output_data_reg[3][4][10]  (.D(\RAM_input_data[3][4] [10]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][4] [10]), .QN());
   DFF_X1 \CNN_output_data_reg[3][4][9]  (.D(\RAM_input_data[3][4] [9]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][4] [9]), .QN());
   DFF_X1 \CNN_output_data_reg[3][4][8]  (.D(\RAM_input_data[3][4] [8]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][4] [8]), .QN());
   DFF_X1 \CNN_output_data_reg[3][4][7]  (.D(\RAM_input_data[3][4] [7]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][4] [7]), .QN());
   DFF_X1 \CNN_output_data_reg[3][4][6]  (.D(\RAM_input_data[3][4] [6]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][4] [6]), .QN());
   DFF_X1 \CNN_output_data_reg[3][4][5]  (.D(\RAM_input_data[3][4] [5]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][4] [5]), .QN());
   DFF_X1 \CNN_output_data_reg[3][4][4]  (.D(\RAM_input_data[3][4] [4]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][4] [4]), .QN());
   DFF_X1 \CNN_output_data_reg[3][4][3]  (.D(\RAM_input_data[3][4] [3]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][4] [3]), .QN());
   DFF_X1 \CNN_output_data_reg[3][4][2]  (.D(\RAM_input_data[3][4] [2]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][4] [2]), .QN());
   DFF_X1 \CNN_output_data_reg[3][4][1]  (.D(\RAM_input_data[3][4] [1]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][4] [1]), .QN());
   DFF_X1 \CNN_output_data_reg[3][4][0]  (.D(\RAM_input_data[3][4] [0]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][4] [0]), .QN());
   DFF_X1 \CNN_output_data_reg[3][3][15]  (.D(\RAM_input_data[3][3] [15]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][3] [15]), .QN());
   DFF_X1 \CNN_output_data_reg[3][3][14]  (.D(\RAM_input_data[3][3] [14]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][3] [14]), .QN());
   DFF_X1 \CNN_output_data_reg[3][3][13]  (.D(\RAM_input_data[3][3] [13]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][3] [13]), .QN());
   DFF_X1 \CNN_output_data_reg[3][3][12]  (.D(\RAM_input_data[3][3] [12]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][3] [12]), .QN());
   DFF_X1 \CNN_output_data_reg[3][3][11]  (.D(\RAM_input_data[3][3] [11]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][3] [11]), .QN());
   DFF_X1 \CNN_output_data_reg[3][3][10]  (.D(\RAM_input_data[3][3] [10]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][3] [10]), .QN());
   DFF_X1 \CNN_output_data_reg[3][3][9]  (.D(\RAM_input_data[3][3] [9]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][3] [9]), .QN());
   DFF_X1 \CNN_output_data_reg[3][3][8]  (.D(\RAM_input_data[3][3] [8]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][3] [8]), .QN());
   DFF_X1 \CNN_output_data_reg[3][3][7]  (.D(\RAM_input_data[3][3] [7]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][3] [7]), .QN());
   DFF_X1 \CNN_output_data_reg[3][3][6]  (.D(\RAM_input_data[3][3] [6]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][3] [6]), .QN());
   DFF_X1 \CNN_output_data_reg[3][3][5]  (.D(\RAM_input_data[3][3] [5]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][3] [5]), .QN());
   DFF_X1 \CNN_output_data_reg[3][3][4]  (.D(\RAM_input_data[3][3] [4]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][3] [4]), .QN());
   DFF_X1 \CNN_output_data_reg[3][3][3]  (.D(\RAM_input_data[3][3] [3]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][3] [3]), .QN());
   DFF_X1 \CNN_output_data_reg[3][3][2]  (.D(\RAM_input_data[3][3] [2]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][3] [2]), .QN());
   DFF_X1 \CNN_output_data_reg[3][3][1]  (.D(\RAM_input_data[3][3] [1]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][3] [1]), .QN());
   DFF_X1 \CNN_output_data_reg[3][3][0]  (.D(\RAM_input_data[3][3] [0]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][3] [0]), .QN());
   DFF_X1 \CNN_output_data_reg[3][2][15]  (.D(\RAM_input_data[3][2] [15]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][2] [15]), .QN());
   DFF_X1 \CNN_output_data_reg[3][2][14]  (.D(\RAM_input_data[3][2] [14]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][2] [14]), .QN());
   DFF_X1 \CNN_output_data_reg[3][2][13]  (.D(\RAM_input_data[3][2] [13]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][2] [13]), .QN());
   DFF_X1 \CNN_output_data_reg[3][2][12]  (.D(\RAM_input_data[3][2] [12]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][2] [12]), .QN());
   DFF_X1 \CNN_output_data_reg[3][2][11]  (.D(\RAM_input_data[3][2] [11]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][2] [11]), .QN());
   DFF_X1 \CNN_output_data_reg[3][2][10]  (.D(\RAM_input_data[3][2] [10]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][2] [10]), .QN());
   DFF_X1 \CNN_output_data_reg[3][2][9]  (.D(\RAM_input_data[3][2] [9]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][2] [9]), .QN());
   DFF_X1 \CNN_output_data_reg[3][2][8]  (.D(\RAM_input_data[3][2] [8]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][2] [8]), .QN());
   DFF_X1 \CNN_output_data_reg[3][2][7]  (.D(\RAM_input_data[3][2] [7]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][2] [7]), .QN());
   DFF_X1 \CNN_output_data_reg[3][2][6]  (.D(\RAM_input_data[3][2] [6]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][2] [6]), .QN());
   DFF_X1 \CNN_output_data_reg[3][2][5]  (.D(\RAM_input_data[3][2] [5]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][2] [5]), .QN());
   DFF_X1 \CNN_output_data_reg[3][2][4]  (.D(\RAM_input_data[3][2] [4]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][2] [4]), .QN());
   DFF_X1 \CNN_output_data_reg[3][2][3]  (.D(\RAM_input_data[3][2] [3]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][2] [3]), .QN());
   DFF_X1 \CNN_output_data_reg[3][2][2]  (.D(\RAM_input_data[3][2] [2]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][2] [2]), .QN());
   DFF_X1 \CNN_output_data_reg[3][2][1]  (.D(\RAM_input_data[3][2] [1]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][2] [1]), .QN());
   DFF_X1 \CNN_output_data_reg[3][2][0]  (.D(\RAM_input_data[3][2] [0]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][2] [0]), .QN());
   DFF_X1 \CNN_output_data_reg[3][1][15]  (.D(\RAM_input_data[3][1] [15]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][1] [15]), .QN());
   DFF_X1 \CNN_output_data_reg[3][1][14]  (.D(\RAM_input_data[3][1] [14]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][1] [14]), .QN());
   DFF_X1 \CNN_output_data_reg[3][1][13]  (.D(\RAM_input_data[3][1] [13]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][1] [13]), .QN());
   DFF_X1 \CNN_output_data_reg[3][1][12]  (.D(\RAM_input_data[3][1] [12]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][1] [12]), .QN());
   DFF_X1 \CNN_output_data_reg[3][1][11]  (.D(\RAM_input_data[3][1] [11]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][1] [11]), .QN());
   DFF_X1 \CNN_output_data_reg[3][1][10]  (.D(\RAM_input_data[3][1] [10]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][1] [10]), .QN());
   DFF_X1 \CNN_output_data_reg[3][1][9]  (.D(\RAM_input_data[3][1] [9]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][1] [9]), .QN());
   DFF_X1 \CNN_output_data_reg[3][1][8]  (.D(\RAM_input_data[3][1] [8]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][1] [8]), .QN());
   DFF_X1 \CNN_output_data_reg[3][1][7]  (.D(\RAM_input_data[3][1] [7]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][1] [7]), .QN());
   DFF_X1 \CNN_output_data_reg[3][1][6]  (.D(\RAM_input_data[3][1] [6]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][1] [6]), .QN());
   DFF_X1 \CNN_output_data_reg[3][1][5]  (.D(\RAM_input_data[3][1] [5]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][1] [5]), .QN());
   DFF_X1 \CNN_output_data_reg[3][1][4]  (.D(\RAM_input_data[3][1] [4]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][1] [4]), .QN());
   DFF_X1 \CNN_output_data_reg[3][1][3]  (.D(\RAM_input_data[3][1] [3]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][1] [3]), .QN());
   DFF_X1 \CNN_output_data_reg[3][1][2]  (.D(\RAM_input_data[3][1] [2]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][1] [2]), .QN());
   DFF_X1 \CNN_output_data_reg[3][1][1]  (.D(\RAM_input_data[3][1] [1]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][1] [1]), .QN());
   DFF_X1 \CNN_output_data_reg[3][1][0]  (.D(\RAM_input_data[3][1] [0]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][1] [0]), .QN());
   DFF_X1 \CNN_output_data_reg[3][0][15]  (.D(\RAM_input_data[3][0] [15]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][0] [15]), .QN());
   DFF_X1 \CNN_output_data_reg[3][0][14]  (.D(\RAM_input_data[3][0] [14]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][0] [14]), .QN());
   DFF_X1 \CNN_output_data_reg[3][0][13]  (.D(\RAM_input_data[3][0] [13]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][0] [13]), .QN());
   DFF_X1 \CNN_output_data_reg[3][0][12]  (.D(\RAM_input_data[3][0] [12]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][0] [12]), .QN());
   DFF_X1 \CNN_output_data_reg[3][0][11]  (.D(\RAM_input_data[3][0] [11]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][0] [11]), .QN());
   DFF_X1 \CNN_output_data_reg[3][0][10]  (.D(\RAM_input_data[3][0] [10]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][0] [10]), .QN());
   DFF_X1 \CNN_output_data_reg[3][0][9]  (.D(\RAM_input_data[3][0] [9]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][0] [9]), .QN());
   DFF_X1 \CNN_output_data_reg[3][0][8]  (.D(\RAM_input_data[3][0] [8]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][0] [8]), .QN());
   DFF_X1 \CNN_output_data_reg[3][0][7]  (.D(\RAM_input_data[3][0] [7]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][0] [7]), .QN());
   DFF_X1 \CNN_output_data_reg[3][0][6]  (.D(\RAM_input_data[3][0] [6]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][0] [6]), .QN());
   DFF_X1 \CNN_output_data_reg[3][0][5]  (.D(\RAM_input_data[3][0] [5]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][0] [5]), .QN());
   DFF_X1 \CNN_output_data_reg[3][0][4]  (.D(\RAM_input_data[3][0] [4]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][0] [4]), .QN());
   DFF_X1 \CNN_output_data_reg[3][0][3]  (.D(\RAM_input_data[3][0] [3]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][0] [3]), .QN());
   DFF_X1 \CNN_output_data_reg[3][0][2]  (.D(\RAM_input_data[3][0] [2]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][0] [2]), .QN());
   DFF_X1 \CNN_output_data_reg[3][0][1]  (.D(\RAM_input_data[3][0] [1]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][0] [1]), .QN());
   DFF_X1 \CNN_output_data_reg[3][0][0]  (.D(\RAM_input_data[3][0] [0]), 
      .CK(n_1_56), .Q(\CNN_output_data[3][0] [0]), .QN());
   DFF_X1 \CNN_output_data_reg[2][4][15]  (.D(\RAM_input_data[2][4] [15]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][4] [15]), .QN());
   DFF_X1 \CNN_output_data_reg[2][4][14]  (.D(\RAM_input_data[2][4] [14]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][4] [14]), .QN());
   DFF_X1 \CNN_output_data_reg[2][4][13]  (.D(\RAM_input_data[2][4] [13]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][4] [13]), .QN());
   DFF_X1 \CNN_output_data_reg[2][4][12]  (.D(\RAM_input_data[2][4] [12]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][4] [12]), .QN());
   DFF_X1 \CNN_output_data_reg[2][4][11]  (.D(\RAM_input_data[2][4] [11]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][4] [11]), .QN());
   DFF_X1 \CNN_output_data_reg[2][4][10]  (.D(\RAM_input_data[2][4] [10]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][4] [10]), .QN());
   DFF_X1 \CNN_output_data_reg[2][4][9]  (.D(\RAM_input_data[2][4] [9]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][4] [9]), .QN());
   DFF_X1 \CNN_output_data_reg[2][4][8]  (.D(\RAM_input_data[2][4] [8]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][4] [8]), .QN());
   DFF_X1 \CNN_output_data_reg[2][4][7]  (.D(\RAM_input_data[2][4] [7]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][4] [7]), .QN());
   DFF_X1 \CNN_output_data_reg[2][4][6]  (.D(\RAM_input_data[2][4] [6]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][4] [6]), .QN());
   DFF_X1 \CNN_output_data_reg[2][4][5]  (.D(\RAM_input_data[2][4] [5]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][4] [5]), .QN());
   DFF_X1 \CNN_output_data_reg[2][4][4]  (.D(\RAM_input_data[2][4] [4]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][4] [4]), .QN());
   DFF_X1 \CNN_output_data_reg[2][4][3]  (.D(\RAM_input_data[2][4] [3]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][4] [3]), .QN());
   DFF_X1 \CNN_output_data_reg[2][4][2]  (.D(\RAM_input_data[2][4] [2]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][4] [2]), .QN());
   DFF_X1 \CNN_output_data_reg[2][4][1]  (.D(\RAM_input_data[2][4] [1]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][4] [1]), .QN());
   DFF_X1 \CNN_output_data_reg[2][4][0]  (.D(\RAM_input_data[2][4] [0]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][4] [0]), .QN());
   DFF_X1 \CNN_output_data_reg[2][3][15]  (.D(\RAM_input_data[2][3] [15]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][3] [15]), .QN());
   DFF_X1 \CNN_output_data_reg[2][3][14]  (.D(\RAM_input_data[2][3] [14]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][3] [14]), .QN());
   DFF_X1 \CNN_output_data_reg[2][3][13]  (.D(\RAM_input_data[2][3] [13]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][3] [13]), .QN());
   DFF_X1 \CNN_output_data_reg[2][3][12]  (.D(\RAM_input_data[2][3] [12]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][3] [12]), .QN());
   DFF_X1 \CNN_output_data_reg[2][3][11]  (.D(\RAM_input_data[2][3] [11]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][3] [11]), .QN());
   DFF_X1 \CNN_output_data_reg[2][3][10]  (.D(\RAM_input_data[2][3] [10]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][3] [10]), .QN());
   DFF_X1 \CNN_output_data_reg[2][3][9]  (.D(\RAM_input_data[2][3] [9]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][3] [9]), .QN());
   DFF_X1 \CNN_output_data_reg[2][3][8]  (.D(\RAM_input_data[2][3] [8]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][3] [8]), .QN());
   DFF_X1 \CNN_output_data_reg[2][3][7]  (.D(\RAM_input_data[2][3] [7]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][3] [7]), .QN());
   DFF_X1 \CNN_output_data_reg[2][3][6]  (.D(\RAM_input_data[2][3] [6]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][3] [6]), .QN());
   DFF_X1 \CNN_output_data_reg[2][3][5]  (.D(\RAM_input_data[2][3] [5]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][3] [5]), .QN());
   DFF_X1 \CNN_output_data_reg[2][3][4]  (.D(\RAM_input_data[2][3] [4]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][3] [4]), .QN());
   DFF_X1 \CNN_output_data_reg[2][3][3]  (.D(\RAM_input_data[2][3] [3]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][3] [3]), .QN());
   DFF_X1 \CNN_output_data_reg[2][3][2]  (.D(\RAM_input_data[2][3] [2]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][3] [2]), .QN());
   DFF_X1 \CNN_output_data_reg[2][3][1]  (.D(\RAM_input_data[2][3] [1]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][3] [1]), .QN());
   DFF_X1 \CNN_output_data_reg[2][3][0]  (.D(\RAM_input_data[2][3] [0]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][3] [0]), .QN());
   DFF_X1 \CNN_output_data_reg[2][2][15]  (.D(\RAM_input_data[2][2] [15]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][2] [15]), .QN());
   DFF_X1 \CNN_output_data_reg[2][2][14]  (.D(\RAM_input_data[2][2] [14]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][2] [14]), .QN());
   DFF_X1 \CNN_output_data_reg[2][2][13]  (.D(\RAM_input_data[2][2] [13]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][2] [13]), .QN());
   DFF_X1 \CNN_output_data_reg[2][2][12]  (.D(\RAM_input_data[2][2] [12]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][2] [12]), .QN());
   DFF_X1 \CNN_output_data_reg[2][2][11]  (.D(\RAM_input_data[2][2] [11]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][2] [11]), .QN());
   DFF_X1 \CNN_output_data_reg[2][2][10]  (.D(\RAM_input_data[2][2] [10]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][2] [10]), .QN());
   DFF_X1 \CNN_output_data_reg[2][2][9]  (.D(\RAM_input_data[2][2] [9]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][2] [9]), .QN());
   DFF_X1 \CNN_output_data_reg[2][2][8]  (.D(\RAM_input_data[2][2] [8]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][2] [8]), .QN());
   DFF_X1 \CNN_output_data_reg[2][2][7]  (.D(\RAM_input_data[2][2] [7]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][2] [7]), .QN());
   DFF_X1 \CNN_output_data_reg[2][2][6]  (.D(\RAM_input_data[2][2] [6]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][2] [6]), .QN());
   DFF_X1 \CNN_output_data_reg[2][2][5]  (.D(\RAM_input_data[2][2] [5]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][2] [5]), .QN());
   DFF_X1 \CNN_output_data_reg[2][2][4]  (.D(\RAM_input_data[2][2] [4]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][2] [4]), .QN());
   DFF_X1 \CNN_output_data_reg[2][2][3]  (.D(\RAM_input_data[2][2] [3]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][2] [3]), .QN());
   DFF_X1 \CNN_output_data_reg[2][2][2]  (.D(\RAM_input_data[2][2] [2]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][2] [2]), .QN());
   DFF_X1 \CNN_output_data_reg[2][2][1]  (.D(\RAM_input_data[2][2] [1]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][2] [1]), .QN());
   DFF_X1 \CNN_output_data_reg[2][2][0]  (.D(\RAM_input_data[2][2] [0]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][2] [0]), .QN());
   DFF_X1 \CNN_output_data_reg[2][1][15]  (.D(\RAM_input_data[2][1] [15]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][1] [15]), .QN());
   DFF_X1 \CNN_output_data_reg[2][1][14]  (.D(\RAM_input_data[2][1] [14]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][1] [14]), .QN());
   DFF_X1 \CNN_output_data_reg[2][1][13]  (.D(\RAM_input_data[2][1] [13]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][1] [13]), .QN());
   DFF_X1 \CNN_output_data_reg[2][1][12]  (.D(\RAM_input_data[2][1] [12]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][1] [12]), .QN());
   DFF_X1 \CNN_output_data_reg[2][1][11]  (.D(\RAM_input_data[2][1] [11]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][1] [11]), .QN());
   DFF_X1 \CNN_output_data_reg[2][1][10]  (.D(\RAM_input_data[2][1] [10]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][1] [10]), .QN());
   DFF_X1 \CNN_output_data_reg[2][1][9]  (.D(\RAM_input_data[2][1] [9]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][1] [9]), .QN());
   DFF_X1 \CNN_output_data_reg[2][1][8]  (.D(\RAM_input_data[2][1] [8]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][1] [8]), .QN());
   DFF_X1 \CNN_output_data_reg[2][1][7]  (.D(\RAM_input_data[2][1] [7]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][1] [7]), .QN());
   DFF_X1 \CNN_output_data_reg[2][1][6]  (.D(\RAM_input_data[2][1] [6]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][1] [6]), .QN());
   DFF_X1 \CNN_output_data_reg[2][1][5]  (.D(\RAM_input_data[2][1] [5]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][1] [5]), .QN());
   DFF_X1 \CNN_output_data_reg[2][1][4]  (.D(\RAM_input_data[2][1] [4]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][1] [4]), .QN());
   DFF_X1 \CNN_output_data_reg[2][1][3]  (.D(\RAM_input_data[2][1] [3]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][1] [3]), .QN());
   DFF_X1 \CNN_output_data_reg[2][1][2]  (.D(\RAM_input_data[2][1] [2]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][1] [2]), .QN());
   DFF_X1 \CNN_output_data_reg[2][1][1]  (.D(\RAM_input_data[2][1] [1]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][1] [1]), .QN());
   DFF_X1 \CNN_output_data_reg[2][1][0]  (.D(\RAM_input_data[2][1] [0]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][1] [0]), .QN());
   DFF_X1 \CNN_output_data_reg[2][0][15]  (.D(\RAM_input_data[2][0] [15]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][0] [15]), .QN());
   DFF_X1 \CNN_output_data_reg[2][0][14]  (.D(\RAM_input_data[2][0] [14]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][0] [14]), .QN());
   DFF_X1 \CNN_output_data_reg[2][0][13]  (.D(\RAM_input_data[2][0] [13]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][0] [13]), .QN());
   DFF_X1 \CNN_output_data_reg[2][0][12]  (.D(\RAM_input_data[2][0] [12]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][0] [12]), .QN());
   DFF_X1 \CNN_output_data_reg[2][0][11]  (.D(\RAM_input_data[2][0] [11]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][0] [11]), .QN());
   DFF_X1 \CNN_output_data_reg[2][0][10]  (.D(\RAM_input_data[2][0] [10]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][0] [10]), .QN());
   DFF_X1 \CNN_output_data_reg[2][0][9]  (.D(\RAM_input_data[2][0] [9]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][0] [9]), .QN());
   DFF_X1 \CNN_output_data_reg[2][0][8]  (.D(\RAM_input_data[2][0] [8]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][0] [8]), .QN());
   DFF_X1 \CNN_output_data_reg[2][0][7]  (.D(\RAM_input_data[2][0] [7]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][0] [7]), .QN());
   DFF_X1 \CNN_output_data_reg[2][0][6]  (.D(\RAM_input_data[2][0] [6]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][0] [6]), .QN());
   DFF_X1 \CNN_output_data_reg[2][0][5]  (.D(\RAM_input_data[2][0] [5]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][0] [5]), .QN());
   DFF_X1 \CNN_output_data_reg[2][0][4]  (.D(\RAM_input_data[2][0] [4]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][0] [4]), .QN());
   DFF_X1 \CNN_output_data_reg[2][0][3]  (.D(\RAM_input_data[2][0] [3]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][0] [3]), .QN());
   DFF_X1 \CNN_output_data_reg[2][0][2]  (.D(\RAM_input_data[2][0] [2]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][0] [2]), .QN());
   DFF_X1 \CNN_output_data_reg[2][0][1]  (.D(\RAM_input_data[2][0] [1]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][0] [1]), .QN());
   DFF_X1 \CNN_output_data_reg[2][0][0]  (.D(\RAM_input_data[2][0] [0]), 
      .CK(n_1_56), .Q(\CNN_output_data[2][0] [0]), .QN());
   DFF_X1 \CNN_output_data_reg[1][4][15]  (.D(\RAM_input_data[1][4] [15]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][4] [15]), .QN());
   DFF_X1 \CNN_output_data_reg[1][4][14]  (.D(\RAM_input_data[1][4] [14]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][4] [14]), .QN());
   DFF_X1 \CNN_output_data_reg[1][4][13]  (.D(\RAM_input_data[1][4] [13]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][4] [13]), .QN());
   DFF_X1 \CNN_output_data_reg[1][4][12]  (.D(\RAM_input_data[1][4] [12]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][4] [12]), .QN());
   DFF_X1 \CNN_output_data_reg[1][4][11]  (.D(\RAM_input_data[1][4] [11]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][4] [11]), .QN());
   DFF_X1 \CNN_output_data_reg[1][4][10]  (.D(\RAM_input_data[1][4] [10]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][4] [10]), .QN());
   DFF_X1 \CNN_output_data_reg[1][4][9]  (.D(\RAM_input_data[1][4] [9]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][4] [9]), .QN());
   DFF_X1 \CNN_output_data_reg[1][4][8]  (.D(\RAM_input_data[1][4] [8]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][4] [8]), .QN());
   DFF_X1 \CNN_output_data_reg[1][4][7]  (.D(\RAM_input_data[1][4] [7]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][4] [7]), .QN());
   DFF_X1 \CNN_output_data_reg[1][4][6]  (.D(\RAM_input_data[1][4] [6]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][4] [6]), .QN());
   DFF_X1 \CNN_output_data_reg[1][4][5]  (.D(\RAM_input_data[1][4] [5]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][4] [5]), .QN());
   DFF_X1 \CNN_output_data_reg[1][4][4]  (.D(\RAM_input_data[1][4] [4]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][4] [4]), .QN());
   DFF_X1 \CNN_output_data_reg[1][4][3]  (.D(\RAM_input_data[1][4] [3]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][4] [3]), .QN());
   DFF_X1 \CNN_output_data_reg[1][4][2]  (.D(\RAM_input_data[1][4] [2]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][4] [2]), .QN());
   DFF_X1 \CNN_output_data_reg[1][4][1]  (.D(\RAM_input_data[1][4] [1]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][4] [1]), .QN());
   DFF_X1 \CNN_output_data_reg[1][4][0]  (.D(\RAM_input_data[1][4] [0]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][4] [0]), .QN());
   DFF_X1 \CNN_output_data_reg[1][3][15]  (.D(\RAM_input_data[1][3] [15]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][3] [15]), .QN());
   DFF_X1 \CNN_output_data_reg[1][3][14]  (.D(\RAM_input_data[1][3] [14]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][3] [14]), .QN());
   DFF_X1 \CNN_output_data_reg[1][3][13]  (.D(\RAM_input_data[1][3] [13]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][3] [13]), .QN());
   DFF_X1 \CNN_output_data_reg[1][3][12]  (.D(\RAM_input_data[1][3] [12]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][3] [12]), .QN());
   DFF_X1 \CNN_output_data_reg[1][3][11]  (.D(\RAM_input_data[1][3] [11]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][3] [11]), .QN());
   DFF_X1 \CNN_output_data_reg[1][3][10]  (.D(\RAM_input_data[1][3] [10]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][3] [10]), .QN());
   DFF_X1 \CNN_output_data_reg[1][3][9]  (.D(\RAM_input_data[1][3] [9]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][3] [9]), .QN());
   DFF_X1 \CNN_output_data_reg[1][3][8]  (.D(\RAM_input_data[1][3] [8]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][3] [8]), .QN());
   DFF_X1 \CNN_output_data_reg[1][3][7]  (.D(\RAM_input_data[1][3] [7]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][3] [7]), .QN());
   DFF_X1 \CNN_output_data_reg[1][3][6]  (.D(\RAM_input_data[1][3] [6]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][3] [6]), .QN());
   DFF_X1 \CNN_output_data_reg[1][3][5]  (.D(\RAM_input_data[1][3] [5]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][3] [5]), .QN());
   DFF_X1 \CNN_output_data_reg[1][3][4]  (.D(\RAM_input_data[1][3] [4]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][3] [4]), .QN());
   DFF_X1 \CNN_output_data_reg[1][3][3]  (.D(\RAM_input_data[1][3] [3]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][3] [3]), .QN());
   DFF_X1 \CNN_output_data_reg[1][3][2]  (.D(\RAM_input_data[1][3] [2]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][3] [2]), .QN());
   DFF_X1 \CNN_output_data_reg[1][3][1]  (.D(\RAM_input_data[1][3] [1]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][3] [1]), .QN());
   DFF_X1 \CNN_output_data_reg[1][3][0]  (.D(\RAM_input_data[1][3] [0]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][3] [0]), .QN());
   DFF_X1 \CNN_output_data_reg[1][2][15]  (.D(\RAM_input_data[1][2] [15]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][2] [15]), .QN());
   DFF_X1 \CNN_output_data_reg[1][2][14]  (.D(\RAM_input_data[1][2] [14]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][2] [14]), .QN());
   DFF_X1 \CNN_output_data_reg[1][2][13]  (.D(\RAM_input_data[1][2] [13]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][2] [13]), .QN());
   DFF_X1 \CNN_output_data_reg[1][2][12]  (.D(\RAM_input_data[1][2] [12]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][2] [12]), .QN());
   DFF_X1 \CNN_output_data_reg[1][2][11]  (.D(\RAM_input_data[1][2] [11]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][2] [11]), .QN());
   DFF_X1 \CNN_output_data_reg[1][2][10]  (.D(\RAM_input_data[1][2] [10]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][2] [10]), .QN());
   DFF_X1 \CNN_output_data_reg[1][2][9]  (.D(\RAM_input_data[1][2] [9]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][2] [9]), .QN());
   DFF_X1 \CNN_output_data_reg[1][2][8]  (.D(\RAM_input_data[1][2] [8]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][2] [8]), .QN());
   DFF_X1 \CNN_output_data_reg[1][2][7]  (.D(\RAM_input_data[1][2] [7]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][2] [7]), .QN());
   DFF_X1 \CNN_output_data_reg[1][2][6]  (.D(\RAM_input_data[1][2] [6]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][2] [6]), .QN());
   DFF_X1 \CNN_output_data_reg[1][2][5]  (.D(\RAM_input_data[1][2] [5]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][2] [5]), .QN());
   DFF_X1 \CNN_output_data_reg[1][2][4]  (.D(\RAM_input_data[1][2] [4]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][2] [4]), .QN());
   DFF_X1 \CNN_output_data_reg[1][2][3]  (.D(\RAM_input_data[1][2] [3]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][2] [3]), .QN());
   DFF_X1 \CNN_output_data_reg[1][2][2]  (.D(\RAM_input_data[1][2] [2]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][2] [2]), .QN());
   DFF_X1 \CNN_output_data_reg[1][2][1]  (.D(\RAM_input_data[1][2] [1]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][2] [1]), .QN());
   DFF_X1 \CNN_output_data_reg[1][2][0]  (.D(\RAM_input_data[1][2] [0]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][2] [0]), .QN());
   DFF_X1 \CNN_output_data_reg[1][1][15]  (.D(\RAM_input_data[1][1] [15]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][1] [15]), .QN());
   DFF_X1 \CNN_output_data_reg[1][1][14]  (.D(\RAM_input_data[1][1] [14]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][1] [14]), .QN());
   DFF_X1 \CNN_output_data_reg[1][1][13]  (.D(\RAM_input_data[1][1] [13]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][1] [13]), .QN());
   DFF_X1 \CNN_output_data_reg[1][1][12]  (.D(\RAM_input_data[1][1] [12]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][1] [12]), .QN());
   DFF_X1 \CNN_output_data_reg[1][1][11]  (.D(\RAM_input_data[1][1] [11]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][1] [11]), .QN());
   DFF_X1 \CNN_output_data_reg[1][1][10]  (.D(\RAM_input_data[1][1] [10]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][1] [10]), .QN());
   DFF_X1 \CNN_output_data_reg[1][1][9]  (.D(\RAM_input_data[1][1] [9]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][1] [9]), .QN());
   DFF_X1 \CNN_output_data_reg[1][1][8]  (.D(\RAM_input_data[1][1] [8]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][1] [8]), .QN());
   DFF_X1 \CNN_output_data_reg[1][1][7]  (.D(\RAM_input_data[1][1] [7]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][1] [7]), .QN());
   DFF_X1 \CNN_output_data_reg[1][1][6]  (.D(\RAM_input_data[1][1] [6]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][1] [6]), .QN());
   DFF_X1 \CNN_output_data_reg[1][1][5]  (.D(\RAM_input_data[1][1] [5]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][1] [5]), .QN());
   DFF_X1 \CNN_output_data_reg[1][1][4]  (.D(\RAM_input_data[1][1] [4]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][1] [4]), .QN());
   DFF_X1 \CNN_output_data_reg[1][1][3]  (.D(\RAM_input_data[1][1] [3]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][1] [3]), .QN());
   DFF_X1 \CNN_output_data_reg[1][1][2]  (.D(\RAM_input_data[1][1] [2]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][1] [2]), .QN());
   DFF_X1 \CNN_output_data_reg[1][1][1]  (.D(\RAM_input_data[1][1] [1]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][1] [1]), .QN());
   DFF_X1 \CNN_output_data_reg[1][1][0]  (.D(\RAM_input_data[1][1] [0]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][1] [0]), .QN());
   DFF_X1 \CNN_output_data_reg[1][0][15]  (.D(\RAM_input_data[1][0] [15]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][0] [15]), .QN());
   DFF_X1 \CNN_output_data_reg[1][0][14]  (.D(\RAM_input_data[1][0] [14]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][0] [14]), .QN());
   DFF_X1 \CNN_output_data_reg[1][0][13]  (.D(\RAM_input_data[1][0] [13]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][0] [13]), .QN());
   DFF_X1 \CNN_output_data_reg[1][0][12]  (.D(\RAM_input_data[1][0] [12]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][0] [12]), .QN());
   DFF_X1 \CNN_output_data_reg[1][0][11]  (.D(\RAM_input_data[1][0] [11]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][0] [11]), .QN());
   DFF_X1 \CNN_output_data_reg[1][0][10]  (.D(\RAM_input_data[1][0] [10]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][0] [10]), .QN());
   DFF_X1 \CNN_output_data_reg[1][0][9]  (.D(\RAM_input_data[1][0] [9]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][0] [9]), .QN());
   DFF_X1 \CNN_output_data_reg[1][0][8]  (.D(\RAM_input_data[1][0] [8]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][0] [8]), .QN());
   DFF_X1 \CNN_output_data_reg[1][0][7]  (.D(\RAM_input_data[1][0] [7]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][0] [7]), .QN());
   DFF_X1 \CNN_output_data_reg[1][0][6]  (.D(\RAM_input_data[1][0] [6]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][0] [6]), .QN());
   DFF_X1 \CNN_output_data_reg[1][0][5]  (.D(\RAM_input_data[1][0] [5]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][0] [5]), .QN());
   DFF_X1 \CNN_output_data_reg[1][0][4]  (.D(\RAM_input_data[1][0] [4]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][0] [4]), .QN());
   DFF_X1 \CNN_output_data_reg[1][0][3]  (.D(\RAM_input_data[1][0] [3]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][0] [3]), .QN());
   DFF_X1 \CNN_output_data_reg[1][0][2]  (.D(\RAM_input_data[1][0] [2]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][0] [2]), .QN());
   DFF_X1 \CNN_output_data_reg[1][0][1]  (.D(\RAM_input_data[1][0] [1]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][0] [1]), .QN());
   DFF_X1 \CNN_output_data_reg[1][0][0]  (.D(\RAM_input_data[1][0] [0]), 
      .CK(n_1_56), .Q(\CNN_output_data[1][0] [0]), .QN());
   DFF_X1 \CNN_output_data_reg[0][4][15]  (.D(\RAM_input_data[0][4] [15]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][4] [15]), .QN());
   DFF_X1 \CNN_output_data_reg[0][4][14]  (.D(\RAM_input_data[0][4] [14]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][4] [14]), .QN());
   DFF_X1 \CNN_output_data_reg[0][4][13]  (.D(\RAM_input_data[0][4] [13]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][4] [13]), .QN());
   DFF_X1 \CNN_output_data_reg[0][4][12]  (.D(\RAM_input_data[0][4] [12]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][4] [12]), .QN());
   DFF_X1 \CNN_output_data_reg[0][4][11]  (.D(\RAM_input_data[0][4] [11]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][4] [11]), .QN());
   DFF_X1 \CNN_output_data_reg[0][4][10]  (.D(\RAM_input_data[0][4] [10]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][4] [10]), .QN());
   DFF_X1 \CNN_output_data_reg[0][4][9]  (.D(\RAM_input_data[0][4] [9]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][4] [9]), .QN());
   DFF_X1 \CNN_output_data_reg[0][4][8]  (.D(\RAM_input_data[0][4] [8]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][4] [8]), .QN());
   DFF_X1 \CNN_output_data_reg[0][4][7]  (.D(\RAM_input_data[0][4] [7]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][4] [7]), .QN());
   DFF_X1 \CNN_output_data_reg[0][4][6]  (.D(\RAM_input_data[0][4] [6]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][4] [6]), .QN());
   DFF_X1 \CNN_output_data_reg[0][4][5]  (.D(\RAM_input_data[0][4] [5]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][4] [5]), .QN());
   DFF_X1 \CNN_output_data_reg[0][4][4]  (.D(\RAM_input_data[0][4] [4]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][4] [4]), .QN());
   DFF_X1 \CNN_output_data_reg[0][4][3]  (.D(\RAM_input_data[0][4] [3]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][4] [3]), .QN());
   DFF_X1 \CNN_output_data_reg[0][4][2]  (.D(\RAM_input_data[0][4] [2]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][4] [2]), .QN());
   DFF_X1 \CNN_output_data_reg[0][4][1]  (.D(\RAM_input_data[0][4] [1]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][4] [1]), .QN());
   DFF_X1 \CNN_output_data_reg[0][4][0]  (.D(\RAM_input_data[0][4] [0]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][4] [0]), .QN());
   DFF_X1 \CNN_output_data_reg[0][3][15]  (.D(\RAM_input_data[0][3] [15]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][3] [15]), .QN());
   DFF_X1 \CNN_output_data_reg[0][3][14]  (.D(\RAM_input_data[0][3] [14]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][3] [14]), .QN());
   DFF_X1 \CNN_output_data_reg[0][3][13]  (.D(\RAM_input_data[0][3] [13]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][3] [13]), .QN());
   DFF_X1 \CNN_output_data_reg[0][3][12]  (.D(\RAM_input_data[0][3] [12]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][3] [12]), .QN());
   DFF_X1 \CNN_output_data_reg[0][3][11]  (.D(\RAM_input_data[0][3] [11]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][3] [11]), .QN());
   DFF_X1 \CNN_output_data_reg[0][3][10]  (.D(\RAM_input_data[0][3] [10]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][3] [10]), .QN());
   DFF_X1 \CNN_output_data_reg[0][3][9]  (.D(\RAM_input_data[0][3] [9]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][3] [9]), .QN());
   DFF_X1 \CNN_output_data_reg[0][3][8]  (.D(\RAM_input_data[0][3] [8]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][3] [8]), .QN());
   DFF_X1 \CNN_output_data_reg[0][3][7]  (.D(\RAM_input_data[0][3] [7]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][3] [7]), .QN());
   DFF_X1 \CNN_output_data_reg[0][3][6]  (.D(\RAM_input_data[0][3] [6]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][3] [6]), .QN());
   DFF_X1 \CNN_output_data_reg[0][3][5]  (.D(\RAM_input_data[0][3] [5]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][3] [5]), .QN());
   DFF_X1 \CNN_output_data_reg[0][3][4]  (.D(\RAM_input_data[0][3] [4]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][3] [4]), .QN());
   DFF_X1 \CNN_output_data_reg[0][3][3]  (.D(\RAM_input_data[0][3] [3]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][3] [3]), .QN());
   DFF_X1 \CNN_output_data_reg[0][3][2]  (.D(\RAM_input_data[0][3] [2]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][3] [2]), .QN());
   DFF_X1 \CNN_output_data_reg[0][3][1]  (.D(\RAM_input_data[0][3] [1]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][3] [1]), .QN());
   DFF_X1 \CNN_output_data_reg[0][3][0]  (.D(\RAM_input_data[0][3] [0]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][3] [0]), .QN());
   DFF_X1 \CNN_output_data_reg[0][2][15]  (.D(\RAM_input_data[0][2] [15]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][2] [15]), .QN());
   DFF_X1 \CNN_output_data_reg[0][2][14]  (.D(\RAM_input_data[0][2] [14]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][2] [14]), .QN());
   DFF_X1 \CNN_output_data_reg[0][2][13]  (.D(\RAM_input_data[0][2] [13]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][2] [13]), .QN());
   DFF_X1 \CNN_output_data_reg[0][2][12]  (.D(\RAM_input_data[0][2] [12]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][2] [12]), .QN());
   DFF_X1 \CNN_output_data_reg[0][2][11]  (.D(\RAM_input_data[0][2] [11]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][2] [11]), .QN());
   DFF_X1 \CNN_output_data_reg[0][2][10]  (.D(\RAM_input_data[0][2] [10]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][2] [10]), .QN());
   DFF_X1 \CNN_output_data_reg[0][2][9]  (.D(\RAM_input_data[0][2] [9]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][2] [9]), .QN());
   DFF_X1 \CNN_output_data_reg[0][2][8]  (.D(\RAM_input_data[0][2] [8]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][2] [8]), .QN());
   DFF_X1 \CNN_output_data_reg[0][2][7]  (.D(\RAM_input_data[0][2] [7]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][2] [7]), .QN());
   DFF_X1 \CNN_output_data_reg[0][2][6]  (.D(\RAM_input_data[0][2] [6]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][2] [6]), .QN());
   DFF_X1 \CNN_output_data_reg[0][2][5]  (.D(\RAM_input_data[0][2] [5]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][2] [5]), .QN());
   DFF_X1 \CNN_output_data_reg[0][2][4]  (.D(\RAM_input_data[0][2] [4]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][2] [4]), .QN());
   DFF_X1 \CNN_output_data_reg[0][2][3]  (.D(\RAM_input_data[0][2] [3]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][2] [3]), .QN());
   DFF_X1 \CNN_output_data_reg[0][2][2]  (.D(\RAM_input_data[0][2] [2]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][2] [2]), .QN());
   DFF_X1 \CNN_output_data_reg[0][2][1]  (.D(\RAM_input_data[0][2] [1]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][2] [1]), .QN());
   DFF_X1 \CNN_output_data_reg[0][2][0]  (.D(\RAM_input_data[0][2] [0]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][2] [0]), .QN());
   DFF_X1 \CNN_output_data_reg[0][1][15]  (.D(\RAM_input_data[0][1] [15]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][1] [15]), .QN());
   DFF_X1 \CNN_output_data_reg[0][1][14]  (.D(\RAM_input_data[0][1] [14]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][1] [14]), .QN());
   DFF_X1 \CNN_output_data_reg[0][1][13]  (.D(\RAM_input_data[0][1] [13]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][1] [13]), .QN());
   DFF_X1 \CNN_output_data_reg[0][1][12]  (.D(\RAM_input_data[0][1] [12]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][1] [12]), .QN());
   DFF_X1 \CNN_output_data_reg[0][1][11]  (.D(\RAM_input_data[0][1] [11]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][1] [11]), .QN());
   DFF_X1 \CNN_output_data_reg[0][1][10]  (.D(\RAM_input_data[0][1] [10]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][1] [10]), .QN());
   DFF_X1 \CNN_output_data_reg[0][1][9]  (.D(\RAM_input_data[0][1] [9]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][1] [9]), .QN());
   DFF_X1 \CNN_output_data_reg[0][1][8]  (.D(\RAM_input_data[0][1] [8]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][1] [8]), .QN());
   DFF_X1 \CNN_output_data_reg[0][1][7]  (.D(\RAM_input_data[0][1] [7]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][1] [7]), .QN());
   DFF_X1 \CNN_output_data_reg[0][1][6]  (.D(\RAM_input_data[0][1] [6]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][1] [6]), .QN());
   DFF_X1 \CNN_output_data_reg[0][1][5]  (.D(\RAM_input_data[0][1] [5]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][1] [5]), .QN());
   DFF_X1 \CNN_output_data_reg[0][1][4]  (.D(\RAM_input_data[0][1] [4]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][1] [4]), .QN());
   DFF_X1 \CNN_output_data_reg[0][1][3]  (.D(\RAM_input_data[0][1] [3]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][1] [3]), .QN());
   DFF_X1 \CNN_output_data_reg[0][1][2]  (.D(\RAM_input_data[0][1] [2]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][1] [2]), .QN());
   DFF_X1 \CNN_output_data_reg[0][1][1]  (.D(\RAM_input_data[0][1] [1]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][1] [1]), .QN());
   DFF_X1 \CNN_output_data_reg[0][1][0]  (.D(\RAM_input_data[0][1] [0]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][1] [0]), .QN());
   DFF_X1 \CNN_output_data_reg[0][0][15]  (.D(\RAM_input_data[0][0] [15]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][0] [15]), .QN());
   DFF_X1 \CNN_output_data_reg[0][0][14]  (.D(\RAM_input_data[0][0] [14]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][0] [14]), .QN());
   DFF_X1 \CNN_output_data_reg[0][0][13]  (.D(\RAM_input_data[0][0] [13]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][0] [13]), .QN());
   DFF_X1 \CNN_output_data_reg[0][0][12]  (.D(\RAM_input_data[0][0] [12]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][0] [12]), .QN());
   DFF_X1 \CNN_output_data_reg[0][0][11]  (.D(\RAM_input_data[0][0] [11]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][0] [11]), .QN());
   DFF_X1 \CNN_output_data_reg[0][0][10]  (.D(\RAM_input_data[0][0] [10]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][0] [10]), .QN());
   DFF_X1 \CNN_output_data_reg[0][0][9]  (.D(\RAM_input_data[0][0] [9]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][0] [9]), .QN());
   DFF_X1 \CNN_output_data_reg[0][0][8]  (.D(\RAM_input_data[0][0] [8]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][0] [8]), .QN());
   DFF_X1 \CNN_output_data_reg[0][0][7]  (.D(\RAM_input_data[0][0] [7]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][0] [7]), .QN());
   DFF_X1 \CNN_output_data_reg[0][0][6]  (.D(\RAM_input_data[0][0] [6]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][0] [6]), .QN());
   DFF_X1 \CNN_output_data_reg[0][0][5]  (.D(\RAM_input_data[0][0] [5]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][0] [5]), .QN());
   DFF_X1 \CNN_output_data_reg[0][0][4]  (.D(\RAM_input_data[0][0] [4]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][0] [4]), .QN());
   DFF_X1 \CNN_output_data_reg[0][0][3]  (.D(\RAM_input_data[0][0] [3]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][0] [3]), .QN());
   DFF_X1 \CNN_output_data_reg[0][0][2]  (.D(\RAM_input_data[0][0] [2]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][0] [2]), .QN());
   DFF_X1 \CNN_output_data_reg[0][0][1]  (.D(\RAM_input_data[0][0] [1]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][0] [1]), .QN());
   DFF_X1 \CNN_output_data_reg[0][0][0]  (.D(\RAM_input_data[0][0] [0]), 
      .CK(n_1_56), .Q(\CNN_output_data[0][0] [0]), .QN());
   CLKGATETST_X1 \clk_gate_CNN_output_data_reg[4][4]_reg  (.CK(clk), .E(n_1_5), 
      .SE(1'b0), .GCK(n_1_56));
   CLKGATETST_X1 clk_gate_biasCounter_reg (.CK(clk), .E(n_1_4), .SE(1'b0), 
      .GCK(n_1_57));
   DFF_X1 \biasCounter_reg[31]  (.D(n_1_3), .CK(n_1_57), .Q(biasCounter[31]), 
      .QN());
   DFF_X1 \biasCounter_reg[2]  (.D(n_1_2), .CK(n_1_57), .Q(biasCounter[2]), 
      .QN());
   DFF_X1 \biasCounter_reg[1]  (.D(n_1_1), .CK(n_1_57), .Q(biasCounter[1]), 
      .QN());
   DFF_X1 \biasCounter_reg[0]  (.D(n_1_0), .CK(n_1_57), .Q(biasCounter[0]), 
      .QN());
   CLKGATETST_X1 clk_gate_inner_address_reg (.CK(clk), .E(n_1_53), .SE(1'b0), 
      .GCK(n_1_58));
   DFF_X1 \inner_address_reg[15]  (.D(n_1_76), .CK(n_1_58), .Q(inner_address[15]), 
      .QN());
   DFF_X1 \inner_address_reg[14]  (.D(n_1_75), .CK(n_1_58), .Q(inner_address[14]), 
      .QN());
   DFF_X1 \inner_address_reg[13]  (.D(n_1_74), .CK(n_1_58), .Q(inner_address[13]), 
      .QN());
   DFF_X1 \inner_address_reg[12]  (.D(n_1_73), .CK(n_1_58), .Q(inner_address[12]), 
      .QN());
   DFF_X1 \inner_address_reg[11]  (.D(n_1_72), .CK(n_1_58), .Q(inner_address[11]), 
      .QN());
   DFF_X1 \inner_address_reg[10]  (.D(n_1_71), .CK(n_1_58), .Q(inner_address[10]), 
      .QN());
   DFF_X1 \inner_address_reg[9]  (.D(n_1_70), .CK(n_1_58), .Q(inner_address[9]), 
      .QN());
   DFF_X1 \inner_address_reg[8]  (.D(n_1_69), .CK(n_1_58), .Q(inner_address[8]), 
      .QN());
   DFF_X1 \inner_address_reg[7]  (.D(n_1_68), .CK(n_1_58), .Q(inner_address[7]), 
      .QN());
   DFF_X1 \inner_address_reg[6]  (.D(n_1_67), .CK(n_1_58), .Q(inner_address[6]), 
      .QN());
   DFF_X1 \inner_address_reg[5]  (.D(n_1_66), .CK(n_1_58), .Q(inner_address[5]), 
      .QN());
   DFF_X1 \inner_address_reg[4]  (.D(n_1_65), .CK(n_1_58), .Q(inner_address[4]), 
      .QN());
   DFF_X1 \inner_address_reg[3]  (.D(n_1_64), .CK(n_1_58), .Q(inner_address[3]), 
      .QN());
   DFF_X1 \inner_address_reg[2]  (.D(n_1_63), .CK(n_1_58), .Q(inner_address[2]), 
      .QN());
   DFF_X1 \inner_address_reg[1]  (.D(n_1_62), .CK(n_1_58), .Q(inner_address[1]), 
      .QN());
   DFF_X1 \inner_address_reg[0]  (.D(n_1_61), .CK(n_1_58), .Q(inner_address[0]), 
      .QN());
   DFF_X1 \RAM_address_reg[15]  (.D(n_1_20), .CK(n_1_59), .Q(n_0), .QN());
   DFF_X1 \RAM_address_reg[14]  (.D(n_1_19), .CK(n_1_59), .Q(n_1), .QN());
   DFF_X1 \RAM_address_reg[13]  (.D(n_1_18), .CK(n_1_59), .Q(n_2), .QN());
   DFF_X1 \RAM_address_reg[12]  (.D(n_1_17), .CK(n_1_59), .Q(n_3), .QN());
   DFF_X1 \RAM_address_reg[11]  (.D(n_1_16), .CK(n_1_59), .Q(n_4), .QN());
   DFF_X1 \RAM_address_reg[10]  (.D(n_1_15), .CK(n_1_59), .Q(n_5), .QN());
   DFF_X1 \RAM_address_reg[9]  (.D(n_1_14), .CK(n_1_59), .Q(n_6), .QN());
   DFF_X1 \RAM_address_reg[8]  (.D(n_1_13), .CK(n_1_59), .Q(n_7), .QN());
   DFF_X1 \RAM_address_reg[7]  (.D(n_1_12), .CK(n_1_59), .Q(n_8), .QN());
   DFF_X1 \RAM_address_reg[6]  (.D(n_1_11), .CK(n_1_59), .Q(n_9), .QN());
   DFF_X1 \RAM_address_reg[5]  (.D(n_1_10), .CK(n_1_59), .Q(n_10), .QN());
   DFF_X1 \RAM_address_reg[4]  (.D(n_1_9), .CK(n_1_59), .Q(n_11), .QN());
   DFF_X1 \RAM_address_reg[3]  (.D(n_1_8), .CK(n_1_59), .Q(n_12), .QN());
   DFF_X1 \RAM_address_reg[2]  (.D(n_1_7), .CK(n_1_59), .Q(n_13), .QN());
   DFF_X1 \RAM_address_reg[1]  (.D(n_1_6), .CK(n_1_59), .Q(n_14), .QN());
   DFF_X1 \RAM_address_reg[0]  (.D(n_1_77), .CK(n_1_59), .Q(n_15), .QN());
   CLKGATETST_X1 clk_gate_RAM_address_reg (.CK(clk), .E(n_1_54), .SE(1'b0), 
      .GCK(n_1_59));
   DFF_X1 FB_bias_or_filter_reg (.D(n_1_60), .CK(clk), .Q(FB_bias_or_filter), 
      .QN());
   MUX2_X1 FB_bias_or_filter_reg_enable_mux_0 (.A(FB_bias_or_filter), .B(n_1_55), 
      .S(n_1_78), .Z(n_1_60));
   DFF_X1 \RAM_address_reg[15]__0  (.D(n_0_16), .CK(n_0_0), .Q(n_0), .QN());
   DFF_X1 \RAM_address_reg[14]__0  (.D(n_0_15), .CK(n_0_0), .Q(n_1), .QN());
   DFF_X1 \RAM_address_reg[13]__0  (.D(n_0_14), .CK(n_0_0), .Q(n_2), .QN());
   DFF_X1 \RAM_address_reg[12]__0  (.D(n_0_13), .CK(n_0_0), .Q(n_3), .QN());
   DFF_X1 \RAM_address_reg[11]__0  (.D(n_0_12), .CK(n_0_0), .Q(n_4), .QN());
   DFF_X1 \RAM_address_reg[10]__0  (.D(n_0_11), .CK(n_0_0), .Q(n_5), .QN());
   DFF_X1 \RAM_address_reg[9]__0  (.D(n_0_10), .CK(n_0_0), .Q(n_6), .QN());
   DFF_X1 \RAM_address_reg[8]__0  (.D(n_0_9), .CK(n_0_0), .Q(n_7), .QN());
   DFF_X1 \RAM_address_reg[7]__0  (.D(n_0_8), .CK(n_0_0), .Q(n_8), .QN());
   DFF_X1 \RAM_address_reg[6]__0  (.D(n_0_7), .CK(n_0_0), .Q(n_9), .QN());
   DFF_X1 \RAM_address_reg[5]__0  (.D(n_0_6), .CK(n_0_0), .Q(n_10), .QN());
   DFF_X1 \RAM_address_reg[4]__0  (.D(n_0_5), .CK(n_0_0), .Q(n_11), .QN());
   DFF_X1 \RAM_address_reg[3]__0  (.D(n_0_4), .CK(n_0_0), .Q(n_12), .QN());
   DFF_X1 \RAM_address_reg[2]__0  (.D(n_0_3), .CK(n_0_0), .Q(n_13), .QN());
   DFF_X1 \RAM_address_reg[1]__0  (.D(n_0_2), .CK(n_0_0), .Q(n_14), .QN());
   DFF_X1 \RAM_address_reg[0]__0  (.D(n_0_1), .CK(n_0_0), .Q(n_15), .QN());
   INV_X1 i_0_0_0 (.A(clk), .ZN(n_0_0));
   NAND2_X1 i_0_1_0 (.A1(read_write_filter_bias[0]), .A2(start), .ZN(n_0_1_0));
   NOR2_X1 i_0_1_1 (.A1(n_0_1_0), .A2(read_write_filter_bias[1]), .ZN(n_0_1_1));
   MUX2_X1 i_0_1_2 (.A(n_0), .B(address[15]), .S(n_0_1_1), .Z(n_0_16));
   MUX2_X1 i_0_1_3 (.A(n_1), .B(address[14]), .S(n_0_1_1), .Z(n_0_15));
   MUX2_X1 i_0_1_4 (.A(n_2), .B(address[13]), .S(n_0_1_1), .Z(n_0_14));
   MUX2_X1 i_0_1_5 (.A(n_3), .B(address[12]), .S(n_0_1_1), .Z(n_0_13));
   MUX2_X1 i_0_1_6 (.A(n_4), .B(address[11]), .S(n_0_1_1), .Z(n_0_12));
   MUX2_X1 i_0_1_7 (.A(n_5), .B(address[10]), .S(n_0_1_1), .Z(n_0_11));
   MUX2_X1 i_0_1_8 (.A(n_6), .B(address[9]), .S(n_0_1_1), .Z(n_0_10));
   MUX2_X1 i_0_1_9 (.A(n_7), .B(address[8]), .S(n_0_1_1), .Z(n_0_9));
   MUX2_X1 i_0_1_10 (.A(n_8), .B(address[7]), .S(n_0_1_1), .Z(n_0_8));
   MUX2_X1 i_0_1_11 (.A(n_9), .B(address[6]), .S(n_0_1_1), .Z(n_0_7));
   MUX2_X1 i_0_1_12 (.A(n_10), .B(address[5]), .S(n_0_1_1), .Z(n_0_6));
   MUX2_X1 i_0_1_13 (.A(n_11), .B(address[4]), .S(n_0_1_1), .Z(n_0_5));
   MUX2_X1 i_0_1_14 (.A(n_12), .B(address[3]), .S(n_0_1_1), .Z(n_0_4));
   MUX2_X1 i_0_1_15 (.A(n_13), .B(address[2]), .S(n_0_1_1), .Z(n_0_3));
   MUX2_X1 i_0_1_16 (.A(n_14), .B(address[1]), .S(n_0_1_1), .Z(n_0_2));
   MUX2_X1 i_0_1_17 (.A(n_15), .B(address[0]), .S(n_0_1_1), .Z(n_0_1));
endmodule

module Filter_Buffer_5x5(read, \input_filter[0][0] , \input_filter[0][1] , 
      \input_filter[0][2] , \input_filter[0][3] , \input_filter[0][4] , 
      \input_filter[1][0] , \input_filter[1][1] , \input_filter[1][2] , 
      \input_filter[1][3] , \input_filter[1][4] , \input_filter[2][0] , 
      \input_filter[2][1] , \input_filter[2][2] , \input_filter[2][3] , 
      \input_filter[2][4] , \input_filter[3][0] , \input_filter[3][1] , 
      \input_filter[3][2] , \input_filter[3][3] , \input_filter[3][4] , 
      \input_filter[4][0] , \input_filter[4][1] , \input_filter[4][2] , 
      \input_filter[4][3] , \input_filter[4][4] , finish, \output_filter[0][0] , 
      \output_filter[0][1] , \output_filter[0][2] , \output_filter[0][3] , 
      \output_filter[0][4] , \output_filter[1][0] , \output_filter[1][1] , 
      \output_filter[1][2] , \output_filter[1][3] , \output_filter[1][4] , 
      \output_filter[2][0] , \output_filter[2][1] , \output_filter[2][2] , 
      \output_filter[2][3] , \output_filter[2][4] , \output_filter[3][0] , 
      \output_filter[3][1] , \output_filter[3][2] , \output_filter[3][3] , 
      \output_filter[3][4] , \output_filter[4][0] , \output_filter[4][1] , 
      \output_filter[4][2] , \output_filter[4][3] , \output_filter[4][4] , 
      index_buffer, index_bias, \input_bias[0] , \input_bias[1] , 
      \input_bias[2] , \input_bias[3] , \input_bias[4] , \input_bias[5] , 
      \input_bias[6] , \input_bias[7] , \input_bias[8] , \input_bias[9] , 
      \input_bias[10] , \input_bias[11] , \input_bias[12] , \input_bias[13] , 
      \input_bias[14] , \input_bias[15] , \input_bias[16] , \input_bias[17] , 
      \input_bias[18] , \input_bias[19] , \input_bias[20] , \input_bias[21] , 
      \input_bias[22] , \input_bias[23] , \input_bias[24] , \input_bias[25] , 
      \input_bias[26] , \input_bias[27] , \input_bias[28] , \input_bias[29] , 
      \input_bias[30] , \input_bias[31] , \input_bias[32] , \input_bias[33] , 
      \input_bias[34] , \input_bias[35] , \input_bias[36] , \input_bias[37] , 
      \input_bias[38] , \input_bias[39] , \input_bias[40] , \input_bias[41] , 
      \input_bias[42] , \input_bias[43] , \input_bias[44] , \input_bias[45] , 
      \input_bias[46] , \input_bias[47] , \input_bias[48] , \input_bias[49] , 
      \input_bias[50] , \input_bias[51] , \input_bias[52] , \input_bias[53] , 
      \input_bias[54] , \input_bias[55] , \input_bias[56] , \input_bias[57] , 
      \input_bias[58] , \input_bias[59] , \input_bias[60] , \input_bias[61] , 
      \input_bias[62] , \input_bias[63] , \input_bias[64] , \input_bias[65] , 
      \input_bias[66] , \input_bias[67] , \input_bias[68] , \input_bias[69] , 
      \input_bias[70] , \input_bias[71] , \input_bias[72] , \input_bias[73] , 
      \input_bias[74] , \input_bias[75] , \input_bias[76] , \input_bias[77] , 
      \input_bias[78] , \input_bias[79] , \input_bias[80] , \input_bias[81] , 
      \input_bias[82] , \input_bias[83] , \input_bias[84] , \input_bias[85] , 
      \input_bias[86] , \input_bias[87] , \input_bias[88] , \input_bias[89] , 
      \input_bias[90] , \input_bias[91] , \input_bias[92] , \input_bias[93] , 
      \input_bias[94] , \input_bias[95] , \input_bias[96] , \input_bias[97] , 
      \input_bias[98] , \input_bias[99] , \input_bias[100] , \input_bias[101] , 
      \input_bias[102] , \input_bias[103] , \input_bias[104] , \input_bias[105] , 
      \input_bias[106] , \input_bias[107] , \input_bias[108] , \input_bias[109] , 
      \input_bias[110] , \input_bias[111] , \input_bias[112] , \input_bias[113] , 
      \input_bias[114] , \input_bias[115] , \input_bias[116] , \input_bias[117] , 
      \input_bias[118] , \input_bias[119] , bias_or_filter, output_bias);
   input read;
   input [15:0]\input_filter[0][0] ;
   input [15:0]\input_filter[0][1] ;
   input [15:0]\input_filter[0][2] ;
   input [15:0]\input_filter[0][3] ;
   input [15:0]\input_filter[0][4] ;
   input [15:0]\input_filter[1][0] ;
   input [15:0]\input_filter[1][1] ;
   input [15:0]\input_filter[1][2] ;
   input [15:0]\input_filter[1][3] ;
   input [15:0]\input_filter[1][4] ;
   input [15:0]\input_filter[2][0] ;
   input [15:0]\input_filter[2][1] ;
   input [15:0]\input_filter[2][2] ;
   input [15:0]\input_filter[2][3] ;
   input [15:0]\input_filter[2][4] ;
   input [15:0]\input_filter[3][0] ;
   input [15:0]\input_filter[3][1] ;
   input [15:0]\input_filter[3][2] ;
   input [15:0]\input_filter[3][3] ;
   input [15:0]\input_filter[3][4] ;
   input [15:0]\input_filter[4][0] ;
   input [15:0]\input_filter[4][1] ;
   input [15:0]\input_filter[4][2] ;
   input [15:0]\input_filter[4][3] ;
   input [15:0]\input_filter[4][4] ;
   output finish;
   output [15:0]\output_filter[0][0] ;
   output [15:0]\output_filter[0][1] ;
   output [15:0]\output_filter[0][2] ;
   output [15:0]\output_filter[0][3] ;
   output [15:0]\output_filter[0][4] ;
   output [15:0]\output_filter[1][0] ;
   output [15:0]\output_filter[1][1] ;
   output [15:0]\output_filter[1][2] ;
   output [15:0]\output_filter[1][3] ;
   output [15:0]\output_filter[1][4] ;
   output [15:0]\output_filter[2][0] ;
   output [15:0]\output_filter[2][1] ;
   output [15:0]\output_filter[2][2] ;
   output [15:0]\output_filter[2][3] ;
   output [15:0]\output_filter[2][4] ;
   output [15:0]\output_filter[3][0] ;
   output [15:0]\output_filter[3][1] ;
   output [15:0]\output_filter[3][2] ;
   output [15:0]\output_filter[3][3] ;
   output [15:0]\output_filter[3][4] ;
   output [15:0]\output_filter[4][0] ;
   output [15:0]\output_filter[4][1] ;
   output [15:0]\output_filter[4][2] ;
   output [15:0]\output_filter[4][3] ;
   output [15:0]\output_filter[4][4] ;
   input [15:0]index_buffer;
   input [15:0]index_bias;
   input [15:0]\input_bias[0] ;
   input [15:0]\input_bias[1] ;
   input [15:0]\input_bias[2] ;
   input [15:0]\input_bias[3] ;
   input [15:0]\input_bias[4] ;
   input [15:0]\input_bias[5] ;
   input [15:0]\input_bias[6] ;
   input [15:0]\input_bias[7] ;
   input [15:0]\input_bias[8] ;
   input [15:0]\input_bias[9] ;
   input [15:0]\input_bias[10] ;
   input [15:0]\input_bias[11] ;
   input [15:0]\input_bias[12] ;
   input [15:0]\input_bias[13] ;
   input [15:0]\input_bias[14] ;
   input [15:0]\input_bias[15] ;
   input [15:0]\input_bias[16] ;
   input [15:0]\input_bias[17] ;
   input [15:0]\input_bias[18] ;
   input [15:0]\input_bias[19] ;
   input [15:0]\input_bias[20] ;
   input [15:0]\input_bias[21] ;
   input [15:0]\input_bias[22] ;
   input [15:0]\input_bias[23] ;
   input [15:0]\input_bias[24] ;
   input [15:0]\input_bias[25] ;
   input [15:0]\input_bias[26] ;
   input [15:0]\input_bias[27] ;
   input [15:0]\input_bias[28] ;
   input [15:0]\input_bias[29] ;
   input [15:0]\input_bias[30] ;
   input [15:0]\input_bias[31] ;
   input [15:0]\input_bias[32] ;
   input [15:0]\input_bias[33] ;
   input [15:0]\input_bias[34] ;
   input [15:0]\input_bias[35] ;
   input [15:0]\input_bias[36] ;
   input [15:0]\input_bias[37] ;
   input [15:0]\input_bias[38] ;
   input [15:0]\input_bias[39] ;
   input [15:0]\input_bias[40] ;
   input [15:0]\input_bias[41] ;
   input [15:0]\input_bias[42] ;
   input [15:0]\input_bias[43] ;
   input [15:0]\input_bias[44] ;
   input [15:0]\input_bias[45] ;
   input [15:0]\input_bias[46] ;
   input [15:0]\input_bias[47] ;
   input [15:0]\input_bias[48] ;
   input [15:0]\input_bias[49] ;
   input [15:0]\input_bias[50] ;
   input [15:0]\input_bias[51] ;
   input [15:0]\input_bias[52] ;
   input [15:0]\input_bias[53] ;
   input [15:0]\input_bias[54] ;
   input [15:0]\input_bias[55] ;
   input [15:0]\input_bias[56] ;
   input [15:0]\input_bias[57] ;
   input [15:0]\input_bias[58] ;
   input [15:0]\input_bias[59] ;
   input [15:0]\input_bias[60] ;
   input [15:0]\input_bias[61] ;
   input [15:0]\input_bias[62] ;
   input [15:0]\input_bias[63] ;
   input [15:0]\input_bias[64] ;
   input [15:0]\input_bias[65] ;
   input [15:0]\input_bias[66] ;
   input [15:0]\input_bias[67] ;
   input [15:0]\input_bias[68] ;
   input [15:0]\input_bias[69] ;
   input [15:0]\input_bias[70] ;
   input [15:0]\input_bias[71] ;
   input [15:0]\input_bias[72] ;
   input [15:0]\input_bias[73] ;
   input [15:0]\input_bias[74] ;
   input [15:0]\input_bias[75] ;
   input [15:0]\input_bias[76] ;
   input [15:0]\input_bias[77] ;
   input [15:0]\input_bias[78] ;
   input [15:0]\input_bias[79] ;
   input [15:0]\input_bias[80] ;
   input [15:0]\input_bias[81] ;
   input [15:0]\input_bias[82] ;
   input [15:0]\input_bias[83] ;
   input [15:0]\input_bias[84] ;
   input [15:0]\input_bias[85] ;
   input [15:0]\input_bias[86] ;
   input [15:0]\input_bias[87] ;
   input [15:0]\input_bias[88] ;
   input [15:0]\input_bias[89] ;
   input [15:0]\input_bias[90] ;
   input [15:0]\input_bias[91] ;
   input [15:0]\input_bias[92] ;
   input [15:0]\input_bias[93] ;
   input [15:0]\input_bias[94] ;
   input [15:0]\input_bias[95] ;
   input [15:0]\input_bias[96] ;
   input [15:0]\input_bias[97] ;
   input [15:0]\input_bias[98] ;
   input [15:0]\input_bias[99] ;
   input [15:0]\input_bias[100] ;
   input [15:0]\input_bias[101] ;
   input [15:0]\input_bias[102] ;
   input [15:0]\input_bias[103] ;
   input [15:0]\input_bias[104] ;
   input [15:0]\input_bias[105] ;
   input [15:0]\input_bias[106] ;
   input [15:0]\input_bias[107] ;
   input [15:0]\input_bias[108] ;
   input [15:0]\input_bias[109] ;
   input [15:0]\input_bias[110] ;
   input [15:0]\input_bias[111] ;
   input [15:0]\input_bias[112] ;
   input [15:0]\input_bias[113] ;
   input [15:0]\input_bias[114] ;
   input [15:0]\input_bias[115] ;
   input [15:0]\input_bias[116] ;
   input [15:0]\input_bias[117] ;
   input [15:0]\input_bias[118] ;
   input [15:0]\input_bias[119] ;
   input bias_or_filter;
   output [15:0]output_bias;

   wire [15:0]\buffer[0][3][3] ;
   wire [15:0]\buffer[1][3][3] ;
   wire [15:0]\buffer[2][3][3] ;
   wire [15:0]\buffer[3][3][3] ;
   wire [15:0]\buffer[4][3][3] ;
   wire [15:0]\buffer[5][3][3] ;
   wire [15:0]\buffer[6][3][3] ;
   wire [15:0]\buffer[7][3][3] ;
   wire [15:0]\buffer[8][3][3] ;
   wire [15:0]\buffer[9][3][3] ;
   wire [15:0]\buffer[10][3][3] ;
   wire [15:0]\buffer[11][3][3] ;
   wire [15:0]\buffer[12][3][3] ;
   wire [15:0]\buffer[13][3][3] ;
   wire [15:0]\buffer[14][3][3] ;
   wire [15:0]\buffer[15][3][3] ;
   wire [15:0]\buffer[0][3][4] ;
   wire [15:0]\buffer[1][3][4] ;
   wire [15:0]\buffer[2][3][4] ;
   wire [15:0]\buffer[12][4][3] ;
   wire [15:0]\buffer[11][4][3] ;
   wire [15:0]\buffer[10][4][3] ;
   wire [15:0]\buffer[9][4][3] ;
   wire [15:0]\buffer[8][4][3] ;
   wire [15:0]\buffer[7][4][3] ;
   wire [15:0]\buffer[6][4][3] ;
   wire [15:0]\buffer[5][4][3] ;
   wire [15:0]\buffer[4][4][3] ;
   wire [15:0]\buffer[3][3][4] ;
   wire [15:0]\buffer[4][3][4] ;
   wire [15:0]\buffer[5][3][4] ;
   wire [15:0]\buffer[0][4][3] ;
   wire [15:0]\buffer[15][4][2] ;
   wire [15:0]\buffer[14][4][2] ;
   wire [15:0]\buffer[13][4][2] ;
   wire [15:0]\buffer[12][4][2] ;
   wire [15:0]\buffer[11][4][2] ;
   wire [15:0]\buffer[10][4][2] ;
   wire [15:0]\buffer[9][4][2] ;
   wire [15:0]\buffer[8][4][2] ;
   wire [15:0]\buffer[7][4][2] ;
   wire [15:0]\buffer[6][4][2] ;
   wire [15:0]\buffer[5][4][2] ;
   wire [15:0]\buffer[4][4][2] ;
   wire [15:0]\buffer[3][4][2] ;
   wire [15:0]\buffer[2][4][2] ;
   wire [15:0]\buffer[1][4][2] ;
   wire [15:0]\buffer[0][4][2] ;
   wire [15:0]\buffer[15][4][1] ;
   wire [15:0]\buffer[14][4][1] ;
   wire [15:0]\buffer[13][4][1] ;
   wire [15:0]\buffer[12][4][1] ;
   wire [15:0]\buffer[11][4][1] ;
   wire [15:0]\buffer[10][4][1] ;
   wire [15:0]\buffer[9][4][1] ;
   wire [15:0]\buffer[8][4][1] ;
   wire [15:0]\buffer[7][4][1] ;
   wire [15:0]\buffer[6][4][1] ;
   wire [15:0]\buffer[5][4][1] ;
   wire [15:0]\buffer[4][4][1] ;
   wire [15:0]\buffer[3][4][1] ;
   wire [15:0]\buffer[2][4][1] ;
   wire [15:0]\buffer[1][4][1] ;
   wire [15:0]\buffer[0][4][1] ;
   wire [15:0]\buffer[15][4][0] ;
   wire [15:0]\buffer[14][4][0] ;
   wire [15:0]\buffer[13][4][0] ;
   wire [15:0]\buffer[12][4][0] ;
   wire [15:0]\buffer[11][4][0] ;
   wire [15:0]\buffer[10][4][0] ;
   wire [15:0]\buffer[9][4][0] ;
   wire [15:0]\buffer[8][4][0] ;
   wire [15:0]\buffer[7][4][0] ;
   wire [15:0]\buffer[6][4][0] ;
   wire [15:0]\buffer[5][4][0] ;
   wire [15:0]\buffer[4][4][0] ;
   wire [15:0]\buffer[3][4][0] ;
   wire [15:0]\buffer[2][4][0] ;
   wire [15:0]\buffer[1][4][0] ;
   wire [15:0]\buffer[0][4][0] ;
   wire [15:0]\buffer[15][3][4] ;
   wire [15:0]\buffer[14][3][4] ;
   wire [15:0]\buffer[13][3][4] ;
   wire [15:0]\buffer[12][3][4] ;
   wire [15:0]\buffer[11][3][4] ;
   wire [15:0]\buffer[10][3][4] ;
   wire [15:0]\buffer[9][3][4] ;
   wire [15:0]\buffer[8][3][4] ;
   wire [15:0]\buffer[7][3][4] ;
   wire [15:0]\buffer[6][3][4] ;
   wire n_53_0;
   wire n_53_1;
   wire n_53_2;
   wire n_53_3;
   wire n_53_4;
   wire n_53_5;
   wire n_53_6;
   wire n_53_7;
   wire n_53_8;
   wire n_53_9;
   wire n_53_10;
   wire n_53_11;
   wire n_53_12;
   wire n_53_13;
   wire n_53_14;
   wire n_53_15;
   wire [15:0]\buffer[1][4][3] ;
   wire [15:0]\buffer[2][4][3] ;
   wire [15:0]\buffer[3][4][3] ;
   wire [15:0]\buffer[13][4][3] ;
   wire [15:0]\buffer[14][4][3] ;
   wire [15:0]\buffer[15][4][3] ;
   wire n_54_6;
   wire [15:0]\buffer[0][4][4] ;
   wire [15:0]\buffer[1][4][4] ;
   wire [15:0]\buffer[2][4][4] ;
   wire [15:0]\buffer[3][4][4] ;
   wire n_54_10;
   wire [15:0]\buffer[4][4][4] ;
   wire n_54_11;
   wire [15:0]\buffer[5][4][4] ;
   wire n_54_12;
   wire [15:0]\buffer[6][4][4] ;
   wire n_54_13;
   wire [15:0]\buffer[7][4][4] ;
   wire n_54_14;
   wire [15:0]\buffer[8][4][4] ;
   wire n_54_15;
   wire [15:0]\buffer[9][4][4] ;
   wire n_54_0;
   wire [15:0]\buffer[10][4][4] ;
   wire n_54_1;
   wire [15:0]\buffer[11][4][4] ;
   wire n_54_2;
   wire [15:0]\buffer[12][4][4] ;
   wire [15:0]\buffer[13][4][4] ;
   wire [15:0]\buffer[14][4][4] ;
   wire [15:0]\buffer[15][4][4] ;
   wire [15:0]\buffer[15][0][0] ;
   wire [15:0]\buffer[2][0][0] ;
   wire [15:0]\buffer[1][0][0] ;
   wire n_54_3;
   wire n_54_4;
   wire n_54_5;
   wire n_54_7;
   wire n_54_8;
   wire n_54_9;
   wire [15:0]\buffer[12][3][2] ;
   wire [15:0]\buffer[11][3][2] ;
   wire [15:0]\buffer[10][3][2] ;
   wire [15:0]\buffer[9][3][2] ;
   wire [15:0]\buffer[8][3][2] ;
   wire [15:0]\buffer[7][3][2] ;
   wire [15:0]\buffer[6][3][2] ;
   wire [15:0]\buffer[5][3][2] ;
   wire [15:0]\buffer[4][3][2] ;
   wire [15:0]\buffer[3][3][2] ;
   wire [15:0]\buffer[2][3][2] ;
   wire [15:0]\buffer[1][3][2] ;
   wire [15:0]\buffer[0][3][2] ;
   wire [15:0]\buffer[15][3][1] ;
   wire [15:0]\buffer[14][3][1] ;
   wire [15:0]\buffer[13][3][1] ;
   wire [15:0]\buffer[12][3][1] ;
   wire [15:0]\buffer[11][3][1] ;
   wire [15:0]\buffer[10][3][1] ;
   wire [15:0]\buffer[9][3][1] ;
   wire [15:0]\buffer[8][3][1] ;
   wire [15:0]\buffer[7][3][1] ;
   wire [15:0]\buffer[6][3][1] ;
   wire [15:0]\buffer[5][3][1] ;
   wire [15:0]\buffer[4][3][1] ;
   wire [15:0]\buffer[3][3][1] ;
   wire [15:0]\buffer[2][3][1] ;
   wire [15:0]\buffer[1][3][1] ;
   wire [15:0]\buffer[0][3][1] ;
   wire [15:0]\buffer[15][3][0] ;
   wire [15:0]\buffer[14][3][0] ;
   wire [15:0]\buffer[13][3][0] ;
   wire [15:0]\buffer[12][3][0] ;
   wire [15:0]\buffer[11][3][0] ;
   wire [15:0]\buffer[10][3][0] ;
   wire [15:0]\buffer[9][3][0] ;
   wire [15:0]\buffer[8][3][0] ;
   wire [15:0]\buffer[7][3][0] ;
   wire [15:0]\buffer[6][3][0] ;
   wire [15:0]\buffer[5][3][0] ;
   wire [15:0]\buffer[4][3][0] ;
   wire [15:0]\buffer[3][3][0] ;
   wire [15:0]\buffer[2][3][0] ;
   wire [15:0]\buffer[1][3][0] ;
   wire [15:0]\buffer[0][3][0] ;
   wire [15:0]\buffer[15][2][4] ;
   wire [15:0]\buffer[14][2][4] ;
   wire [15:0]\buffer[13][2][4] ;
   wire [15:0]\buffer[12][2][4] ;
   wire [15:0]\buffer[11][2][4] ;
   wire [15:0]\buffer[10][2][4] ;
   wire [15:0]\buffer[9][2][4] ;
   wire [15:0]\buffer[8][2][4] ;
   wire [15:0]\buffer[7][2][4] ;
   wire [15:0]\buffer[6][2][4] ;
   wire [15:0]\buffer[5][2][4] ;
   wire [15:0]\buffer[4][2][4] ;
   wire [15:0]\buffer[3][2][4] ;
   wire [15:0]\buffer[2][2][4] ;
   wire [15:0]\buffer[1][2][4] ;
   wire [15:0]\buffer[0][2][4] ;
   wire [15:0]\buffer[15][2][3] ;
   wire [15:0]\buffer[14][2][3] ;
   wire [15:0]\buffer[13][2][3] ;
   wire [15:0]\buffer[12][2][3] ;
   wire [15:0]\buffer[11][2][3] ;
   wire [15:0]\buffer[10][2][3] ;
   wire [15:0]\buffer[9][2][3] ;
   wire [15:0]\buffer[8][2][3] ;
   wire [15:0]\buffer[7][2][3] ;
   wire [15:0]\buffer[6][2][3] ;
   wire [15:0]\buffer[5][2][3] ;
   wire [15:0]\buffer[4][2][3] ;
   wire [15:0]\buffer[3][2][3] ;
   wire [15:0]\buffer[2][2][3] ;
   wire [15:0]\buffer[1][2][3] ;
   wire [15:0]\buffer[0][2][3] ;
   wire [15:0]\buffer[15][2][2] ;
   wire [15:0]\buffer[14][2][2] ;
   wire [15:0]\buffer[13][2][2] ;
   wire [15:0]\buffer[12][2][2] ;
   wire [15:0]\buffer[11][2][2] ;
   wire [15:0]\buffer[10][2][2] ;
   wire [15:0]\buffer[9][2][2] ;
   wire [15:0]\buffer[8][2][2] ;
   wire [15:0]\buffer[7][2][2] ;
   wire [15:0]\buffer[6][2][2] ;
   wire [15:0]\buffer[5][2][2] ;
   wire [15:0]\buffer[4][2][2] ;
   wire [15:0]\buffer[3][2][2] ;
   wire [15:0]\buffer[2][2][2] ;
   wire [15:0]\buffer[1][2][2] ;
   wire [15:0]\buffer[0][2][2] ;
   wire [15:0]\buffer[0][0][0] ;
   wire [15:0]\buffer[13][3][2] ;
   wire [15:0]\buffer[14][3][2] ;
   wire [15:0]\buffer[15][3][2] ;
   wire n_55_0;
   wire n_55_1;
   wire n_55_2;
   wire n_55_3;
   wire n_55_4;
   wire n_55_5;
   wire n_55_6;
   wire n_55_7;
   wire n_55_8;
   wire n_55_9;
   wire n_55_10;
   wire n_55_11;
   wire n_55_12;
   wire n_55_13;
   wire n_55_14;
   wire n_55_15;
   wire [15:0]\buffer[3][0][0] ;
   wire [15:0]\buffer[4][0][0] ;
   wire [15:0]\buffer[5][0][0] ;
   wire [15:0]\buffer[6][0][0] ;
   wire [15:0]\buffer[7][0][0] ;
   wire [15:0]\buffer[8][0][0] ;
   wire [15:0]\buffer[9][0][0] ;
   wire [15:0]\buffer[10][0][0] ;
   wire [15:0]\buffer[11][0][0] ;
   wire [15:0]\buffer[12][0][0] ;
   wire [15:0]\buffer[13][0][0] ;
   wire [15:0]\buffer[14][0][0] ;
   wire [15:0]\buffer[0][0][1] ;
   wire [15:0]\buffer[1][0][1] ;
   wire [15:0]\buffer[2][0][1] ;
   wire [15:0]\buffer[3][0][1] ;
   wire [15:0]\buffer[4][0][1] ;
   wire [15:0]\buffer[5][0][1] ;
   wire [15:0]\buffer[6][0][1] ;
   wire [15:0]\buffer[7][0][1] ;
   wire [15:0]\buffer[8][0][1] ;
   wire [15:0]\buffer[9][0][1] ;
   wire [15:0]\buffer[10][0][1] ;
   wire [15:0]\buffer[11][0][1] ;
   wire [15:0]\buffer[12][0][1] ;
   wire [15:0]\buffer[13][0][1] ;
   wire [15:0]\buffer[14][0][1] ;
   wire [15:0]\buffer[15][0][1] ;
   wire [15:0]\buffer[6][0][2] ;
   wire [15:0]\buffer[15][0][2] ;
   wire [15:0]\buffer[1][0][3] ;
   wire [15:0]\buffer[2][0][3] ;
   wire [15:0]\buffer[3][0][3] ;
   wire [15:0]\buffer[10][1][4] ;
   wire [15:0]\buffer[9][1][4] ;
   wire [15:0]\buffer[8][1][4] ;
   wire [15:0]\buffer[7][1][4] ;
   wire [15:0]\buffer[6][1][4] ;
   wire [15:0]\buffer[5][1][4] ;
   wire [15:0]\buffer[4][1][4] ;
   wire [15:0]\buffer[3][1][4] ;
   wire [15:0]\buffer[2][1][4] ;
   wire [15:0]\buffer[1][1][4] ;
   wire [15:0]\buffer[4][0][3] ;
   wire [15:0]\buffer[5][0][3] ;
   wire [15:0]\buffer[6][0][3] ;
   wire [15:0]\buffer[7][0][3] ;
   wire [15:0]\buffer[8][0][3] ;
   wire [15:0]\buffer[9][0][3] ;
   wire [15:0]\buffer[10][0][3] ;
   wire [15:0]\buffer[11][0][3] ;
   wire [15:0]\buffer[12][0][3] ;
   wire [15:0]\buffer[13][0][3] ;
   wire [15:0]\buffer[14][0][3] ;
   wire [15:0]\buffer[15][0][3] ;
   wire [15:0]\buffer[0][1][0] ;
   wire [15:0]\buffer[1][1][0] ;
   wire [15:0]\buffer[2][1][0] ;
   wire [15:0]\buffer[3][1][0] ;
   wire [15:0]\buffer[4][1][0] ;
   wire [15:0]\buffer[5][1][0] ;
   wire [15:0]\buffer[6][1][0] ;
   wire [15:0]\buffer[7][1][0] ;
   wire [15:0]\buffer[8][1][0] ;
   wire [15:0]\buffer[9][1][0] ;
   wire [15:0]\buffer[10][1][0] ;
   wire [15:0]\buffer[11][1][0] ;
   wire [15:0]\buffer[8][1][2] ;
   wire [15:0]\buffer[7][1][2] ;
   wire [15:0]\buffer[6][1][2] ;
   wire [15:0]\buffer[5][1][2] ;
   wire [15:0]\buffer[4][1][2] ;
   wire [15:0]\buffer[3][1][2] ;
   wire [15:0]\buffer[2][1][2] ;
   wire [15:0]\buffer[1][1][2] ;
   wire [15:0]\buffer[12][1][0] ;
   wire [15:0]\buffer[15][1][1] ;
   wire [15:0]\buffer[14][1][1] ;
   wire [15:0]\buffer[13][1][1] ;
   wire [15:0]\buffer[12][1][1] ;
   wire [15:0]\buffer[11][1][1] ;
   wire [15:0]\buffer[10][1][1] ;
   wire [15:0]\buffer[9][1][1] ;
   wire [15:0]\buffer[8][1][1] ;
   wire [15:0]\buffer[7][1][1] ;
   wire [15:0]\buffer[6][1][1] ;
   wire [15:0]\buffer[5][1][1] ;
   wire [15:0]\buffer[4][1][1] ;
   wire [15:0]\buffer[3][1][1] ;
   wire [15:0]\buffer[2][1][1] ;
   wire [15:0]\buffer[1][1][1] ;
   wire [15:0]\buffer[0][1][1] ;
   wire [15:0]\buffer[15][1][0] ;
   wire [15:0]\buffer[14][1][0] ;
   wire [15:0]\buffer[13][1][0] ;
   wire n_56_0;
   wire n_56_1;
   wire n_56_2;
   wire n_56_3;
   wire n_56_4;
   wire n_56_5;
   wire n_56_6;
   wire n_56_7;
   wire n_56_8;
   wire n_56_9;
   wire n_56_10;
   wire n_56_11;
   wire n_56_12;
   wire n_56_13;
   wire n_56_14;
   wire n_56_15;
   wire [15:0]\buffer[0][1][2] ;
   wire [15:0]\buffer[9][1][2] ;
   wire [15:0]\buffer[10][1][2] ;
   wire [15:0]\buffer[11][1][2] ;
   wire [15:0]\buffer[12][1][2] ;
   wire [15:0]\buffer[13][1][2] ;
   wire [15:0]\buffer[14][1][2] ;
   wire [15:0]\buffer[15][1][2] ;
   wire n_57_8;
   wire [15:0]\buffer[4][0][4] ;
   wire n_57_9;
   wire [15:0]\buffer[3][0][4] ;
   wire n_57_10;
   wire [15:0]\buffer[2][0][4] ;
   wire n_57_11;
   wire [15:0]\buffer[1][0][4] ;
   wire [15:0]\buffer[0][0][4] ;
   wire [15:0]\buffer[15][0][4] ;
   wire [15:0]\buffer[14][0][4] ;
   wire [15:0]\buffer[13][0][4] ;
   wire [15:0]\buffer[12][0][4] ;
   wire [15:0]\buffer[11][0][4] ;
   wire [15:0]\buffer[10][0][4] ;
   wire [15:0]\buffer[9][0][4] ;
   wire n_57_0;
   wire [15:0]\buffer[8][0][4] ;
   wire n_57_1;
   wire [15:0]\buffer[7][0][4] ;
   wire n_57_2;
   wire [15:0]\buffer[6][0][4] ;
   wire n_57_3;
   wire [15:0]\buffer[5][0][4] ;
   wire n_57_4;
   wire n_57_5;
   wire n_57_6;
   wire n_57_7;
   wire n_57_12;
   wire n_57_13;
   wire n_57_14;
   wire n_57_15;
   wire [15:0]\buffer[0][1][3] ;
   wire [15:0]\buffer[1][1][3] ;
   wire [15:0]\buffer[2][1][3] ;
   wire [15:0]\buffer[3][1][3] ;
   wire [15:0]\buffer[4][1][3] ;
   wire [15:0]\buffer[5][1][3] ;
   wire n_58_6;
   wire [15:0]\buffer[6][1][3] ;
   wire [15:0]\buffer[7][1][3] ;
   wire [15:0]\buffer[8][1][3] ;
   wire [15:0]\buffer[9][1][3] ;
   wire [15:0]\buffer[10][1][3] ;
   wire [15:0]\buffer[11][1][3] ;
   wire [15:0]\buffer[12][1][3] ;
   wire [15:0]\buffer[13][1][3] ;
   wire [15:0]\buffer[14][1][3] ;
   wire n_58_15;
   wire [15:0]\buffer[15][1][3] ;
   wire [15:0]\buffer[5][0][2] ;
   wire [15:0]\buffer[4][0][2] ;
   wire [15:0]\buffer[3][0][2] ;
   wire [15:0]\buffer[2][0][2] ;
   wire [15:0]\buffer[0][0][3] ;
   wire [15:0]\buffer[1][0][2] ;
   wire [15:0]\buffer[14][0][2] ;
   wire [15:0]\buffer[13][0][2] ;
   wire [15:0]\buffer[12][0][2] ;
   wire [15:0]\buffer[11][0][2] ;
   wire [15:0]\buffer[10][0][2] ;
   wire [15:0]\buffer[9][0][2] ;
   wire [15:0]\buffer[8][0][2] ;
   wire [15:0]\buffer[7][0][2] ;
   wire [15:0]\buffer[0][0][2] ;
   wire n_58_0;
   wire n_58_1;
   wire n_58_2;
   wire n_58_3;
   wire n_58_4;
   wire n_58_5;
   wire n_58_7;
   wire n_58_8;
   wire n_58_9;
   wire n_58_10;
   wire n_58_11;
   wire n_58_12;
   wire n_58_13;
   wire n_58_14;
   wire [15:0]\buffer[0][1][4] ;
   wire [15:0]\buffer[11][1][4] ;
   wire [15:0]\buffer[12][1][4] ;
   wire [15:0]\buffer[13][1][4] ;
   wire [15:0]\buffer[14][1][4] ;
   wire [15:0]\buffer[15][1][4] ;
   wire [15:0]\buffer[0][2][0] ;
   wire [15:0]\buffer[1][2][0] ;
   wire [15:0]\buffer[2][2][0] ;
   wire [15:0]\buffer[3][2][0] ;
   wire [15:0]\buffer[4][2][0] ;
   wire [15:0]\buffer[5][2][0] ;
   wire [15:0]\buffer[6][2][0] ;
   wire [15:0]\buffer[7][2][0] ;
   wire [15:0]\buffer[8][2][0] ;
   wire [15:0]\buffer[9][2][0] ;
   wire [15:0]\buffer[10][2][0] ;
   wire [15:0]\buffer[11][2][0] ;
   wire [15:0]\buffer[12][2][0] ;
   wire [15:0]\buffer[13][2][0] ;
   wire [15:0]\buffer[14][2][0] ;
   wire [15:0]\buffer[15][2][0] ;
   wire [15:0]\buffer[12][2][1] ;
   wire [15:0]\buffer[0][2][1] ;
   wire [15:0]\buffer[1][2][1] ;
   wire [15:0]\buffer[2][2][1] ;
   wire [15:0]\buffer[3][2][1] ;
   wire [15:0]\buffer[4][2][1] ;
   wire [15:0]\buffer[5][2][1] ;
   wire [15:0]\buffer[6][2][1] ;
   wire [15:0]\buffer[7][2][1] ;
   wire [15:0]\buffer[8][2][1] ;
   wire [15:0]\buffer[9][2][1] ;
   wire [15:0]\buffer[10][2][1] ;
   wire [15:0]\buffer[11][2][1] ;
   wire [15:0]\buffer[13][2][1] ;
   wire [15:0]\buffer[14][2][1] ;
   wire [15:0]\buffer[15][2][1] ;
   wire n_59_0;
   wire n_59_1;
   wire n_59_2;
   wire n_59_3;
   wire n_59_4;
   wire n_59_5;
   wire n_59_7;
   wire n_59_8;
   wire n_59_9;
   wire n_59_10;
   wire n_59_11;
   wire n_59_12;
   wire n_59_13;
   wire n_59_14;
   wire n_59_15;
   wire n_59_6;
   wire n_1_0_0;
   wire n_1_0_1;
   wire n_1_0_2;
   wire n_1_0_3;
   wire n_1_0_4;
   wire n_1_0_5;
   wire n_1_0_6;
   wire n_1_0_7;
   wire n_1_0_8;
   wire n_1_0_9;
   wire n_1_0_10;
   wire n_1_0_11;
   wire n_1_0_12;
   wire n_1_0_13;
   wire n_1_0_14;
   wire n_2_44_0;
   wire n_2_44_1;
   wire n_2_44_2;
   wire n_2_44_3;
   wire n_2_44_4;
   wire n_2_44_5;
   wire n_2_44_6;
   wire n_2_44_7;
   wire n_2_44_8;
   wire n_2_44_9;
   wire n_2_44_10;
   wire n_2_44_11;
   wire n_2_44_12;
   wire n_2_44_13;
   wire n_2_44_14;
   wire n_2_44_15;
   wire n_2_44_16;
   wire n_2_44_17;
   wire n_2_44_18;
   wire n_2_44_19;
   wire n_2_44_20;
   wire n_2_44_21;
   wire n_2_44_22;
   wire n_2_44_23;
   wire n_2_44_24;
   wire n_2_44_25;
   wire n_2_44_26;
   wire n_2_44_27;
   wire n_2_44_28;
   wire n_2_44_29;
   wire n_2_44_30;
   wire n_2_44_31;
   wire n_2_44_32;
   wire n_2_44_33;
   wire n_2_44_34;
   wire n_2_44_35;
   wire n_2_44_36;
   wire n_2_44_37;
   wire n_2_44_38;
   wire n_2_44_39;
   wire n_2_44_40;
   wire n_2_44_41;
   wire n_2_44_42;
   wire n_2_44_43;
   wire n_2_44_44;
   wire n_2_44_45;
   wire n_2_44_46;
   wire n_2_44_47;
   wire n_2_44_48;
   wire n_2_44_49;
   wire n_2_44_50;
   wire n_2_44_51;
   wire n_2_44_52;
   wire n_2_44_53;
   wire n_2_44_54;
   wire n_2_44_55;
   wire n_2_44_56;
   wire n_2_44_57;
   wire n_2_44_58;
   wire n_2_44_59;
   wire n_2_44_60;
   wire n_2_44_61;
   wire n_2_44_62;
   wire n_2_44_63;
   wire n_2_44_64;
   wire n_2_44_65;
   wire n_2_44_66;
   wire n_2_44_67;
   wire n_2_44_68;
   wire n_2_44_69;
   wire n_2_44_70;
   wire n_2_44_71;
   wire n_2_44_72;
   wire n_2_44_73;
   wire n_2_44_74;
   wire n_2_44_75;
   wire n_2_44_76;
   wire n_2_44_77;
   wire n_2_44_78;
   wire n_2_44_79;
   wire n_2_44_80;
   wire n_2_44_81;
   wire n_2_44_82;
   wire n_2_44_83;
   wire n_2_44_84;
   wire n_2_44_85;
   wire n_2_44_86;
   wire n_2_44_87;
   wire n_2_44_88;
   wire n_2_44_89;
   wire n_2_44_90;
   wire n_2_44_91;
   wire n_2_44_92;
   wire n_2_44_93;
   wire n_2_44_94;
   wire n_2_44_95;
   wire n_2_44_96;
   wire n_2_44_97;
   wire n_2_44_98;
   wire n_2_44_99;
   wire n_2_44_100;
   wire n_2_44_101;
   wire n_2_44_102;
   wire n_2_44_103;
   wire n_2_44_104;
   wire n_2_44_105;
   wire n_2_44_106;
   wire n_2_44_107;
   wire n_2_44_108;
   wire n_2_44_109;
   wire n_2_44_110;
   wire n_2_44_111;
   wire n_2_44_112;
   wire n_2_44_113;
   wire n_2_44_114;
   wire n_2_44_115;
   wire n_2_44_116;
   wire n_2_44_117;
   wire n_2_44_118;
   wire n_2_44_119;
   wire n_2_44_120;
   wire n_2_44_121;
   wire n_2_44_122;
   wire n_2_44_123;
   wire n_2_44_124;
   wire n_2_44_125;
   wire n_2_44_126;
   wire n_2_44_127;
   wire n_2_44_128;
   wire n_2_44_129;
   wire n_2_44_130;
   wire n_2_44_131;
   wire n_2_44_132;
   wire n_2_44_133;
   wire n_2_44_134;
   wire n_2_44_135;
   wire n_2_44_136;
   wire n_2_44_137;
   wire n_2_44_138;
   wire n_2_44_139;
   wire n_2_44_140;
   wire n_2_44_141;
   wire n_2_44_142;
   wire n_2_44_143;
   wire n_2_44_144;
   wire n_3_43_0;
   wire n_3_43_1;
   wire n_3_43_2;
   wire n_3_43_3;
   wire n_3_43_4;
   wire n_3_43_5;
   wire n_3_43_6;
   wire n_3_43_7;
   wire n_3_43_8;
   wire n_3_43_9;
   wire n_3_43_10;
   wire n_3_43_11;
   wire n_3_43_12;
   wire n_3_43_13;
   wire n_3_43_14;
   wire n_3_43_15;
   wire n_3_43_16;
   wire n_3_43_17;
   wire n_3_43_18;
   wire n_3_43_19;
   wire n_3_43_20;
   wire n_3_43_21;
   wire n_3_43_22;
   wire n_3_43_23;
   wire n_3_43_24;
   wire n_3_43_25;
   wire n_3_43_26;
   wire n_3_43_27;
   wire n_3_43_28;
   wire n_3_43_29;
   wire n_3_43_30;
   wire n_3_43_31;
   wire n_3_43_32;
   wire n_3_43_33;
   wire n_3_43_34;
   wire n_3_43_35;
   wire n_3_43_36;
   wire n_3_43_37;
   wire n_3_43_38;
   wire n_3_43_39;
   wire n_3_43_40;
   wire n_3_43_41;
   wire n_3_43_42;
   wire n_3_43_43;
   wire n_3_43_44;
   wire n_3_43_45;
   wire n_3_43_46;
   wire n_3_43_47;
   wire n_3_43_48;
   wire n_3_43_49;
   wire n_3_43_50;
   wire n_3_43_51;
   wire n_3_43_52;
   wire n_3_43_53;
   wire n_3_43_54;
   wire n_3_43_55;
   wire n_3_43_56;
   wire n_3_43_57;
   wire n_3_43_58;
   wire n_3_43_59;
   wire n_3_43_60;
   wire n_3_43_61;
   wire n_3_43_62;
   wire n_3_43_63;
   wire n_3_43_64;
   wire n_3_43_65;
   wire n_3_43_66;
   wire n_3_43_67;
   wire n_3_43_68;
   wire n_3_43_69;
   wire n_3_43_70;
   wire n_3_43_71;
   wire n_3_43_72;
   wire n_3_43_73;
   wire n_3_43_74;
   wire n_3_43_75;
   wire n_3_43_76;
   wire n_3_43_77;
   wire n_3_43_78;
   wire n_3_43_79;
   wire n_3_43_80;
   wire n_3_43_81;
   wire n_3_43_82;
   wire n_3_43_83;
   wire n_3_43_84;
   wire n_3_43_85;
   wire n_3_43_86;
   wire n_3_43_87;
   wire n_3_43_88;
   wire n_3_43_89;
   wire n_3_43_90;
   wire n_3_43_91;
   wire n_3_43_92;
   wire n_3_43_93;
   wire n_3_43_94;
   wire n_3_43_95;
   wire n_3_43_96;
   wire n_3_43_97;
   wire n_3_43_98;
   wire n_3_43_99;
   wire n_3_43_100;
   wire n_3_43_101;
   wire n_3_43_102;
   wire n_3_43_103;
   wire n_3_43_104;
   wire n_3_43_105;
   wire n_3_43_106;
   wire n_3_43_107;
   wire n_3_43_108;
   wire n_3_43_109;
   wire n_3_43_110;
   wire n_3_43_111;
   wire n_3_43_112;
   wire n_3_43_113;
   wire n_3_43_114;
   wire n_3_43_115;
   wire n_3_43_116;
   wire n_3_43_117;
   wire n_3_43_118;
   wire n_3_43_119;
   wire n_3_43_120;
   wire n_3_43_121;
   wire n_3_43_122;
   wire n_3_43_123;
   wire n_3_43_124;
   wire n_3_43_125;
   wire n_3_43_126;
   wire n_3_43_127;
   wire n_3_43_128;
   wire n_3_43_129;
   wire n_3_43_130;
   wire n_3_43_131;
   wire n_3_43_132;
   wire n_3_43_133;
   wire n_3_43_134;
   wire n_3_43_135;
   wire n_3_43_136;
   wire n_3_43_137;
   wire n_3_43_138;
   wire n_3_43_139;
   wire n_3_43_140;
   wire n_3_43_141;
   wire n_3_43_142;
   wire n_3_43_143;
   wire n_3_43_144;
   wire n_4_42_0;
   wire n_4_42_1;
   wire n_4_42_2;
   wire n_4_42_3;
   wire n_4_42_4;
   wire n_4_42_5;
   wire n_4_42_6;
   wire n_4_42_7;
   wire n_4_42_8;
   wire n_4_42_9;
   wire n_4_42_10;
   wire n_4_42_11;
   wire n_4_42_12;
   wire n_4_42_13;
   wire n_4_42_14;
   wire n_4_42_15;
   wire n_4_42_16;
   wire n_4_42_17;
   wire n_4_42_18;
   wire n_4_42_19;
   wire n_4_42_20;
   wire n_4_42_21;
   wire n_4_42_22;
   wire n_4_42_23;
   wire n_4_42_24;
   wire n_4_42_25;
   wire n_4_42_26;
   wire n_4_42_27;
   wire n_4_42_28;
   wire n_4_42_29;
   wire n_4_42_30;
   wire n_4_42_31;
   wire n_4_42_32;
   wire n_4_42_33;
   wire n_4_42_34;
   wire n_4_42_35;
   wire n_4_42_36;
   wire n_4_42_37;
   wire n_4_42_38;
   wire n_4_42_39;
   wire n_4_42_40;
   wire n_4_42_41;
   wire n_4_42_42;
   wire n_4_42_43;
   wire n_4_42_44;
   wire n_4_42_45;
   wire n_4_42_46;
   wire n_4_42_47;
   wire n_4_42_48;
   wire n_4_42_49;
   wire n_4_42_50;
   wire n_4_42_51;
   wire n_4_42_52;
   wire n_4_42_53;
   wire n_4_42_54;
   wire n_4_42_55;
   wire n_4_42_56;
   wire n_4_42_57;
   wire n_4_42_58;
   wire n_4_42_59;
   wire n_4_42_60;
   wire n_4_42_61;
   wire n_4_42_62;
   wire n_4_42_63;
   wire n_4_42_64;
   wire n_4_42_65;
   wire n_4_42_66;
   wire n_4_42_67;
   wire n_4_42_68;
   wire n_4_42_69;
   wire n_4_42_70;
   wire n_4_42_71;
   wire n_4_42_72;
   wire n_4_42_73;
   wire n_4_42_74;
   wire n_4_42_75;
   wire n_4_42_76;
   wire n_4_42_77;
   wire n_4_42_78;
   wire n_4_42_79;
   wire n_4_42_80;
   wire n_4_42_81;
   wire n_4_42_82;
   wire n_4_42_83;
   wire n_4_42_84;
   wire n_4_42_85;
   wire n_4_42_86;
   wire n_4_42_87;
   wire n_4_42_88;
   wire n_4_42_89;
   wire n_4_42_90;
   wire n_4_42_91;
   wire n_4_42_92;
   wire n_4_42_93;
   wire n_4_42_94;
   wire n_4_42_95;
   wire n_4_42_96;
   wire n_4_42_97;
   wire n_4_42_98;
   wire n_4_42_99;
   wire n_4_42_100;
   wire n_4_42_101;
   wire n_4_42_102;
   wire n_4_42_103;
   wire n_4_42_104;
   wire n_4_42_105;
   wire n_4_42_106;
   wire n_4_42_107;
   wire n_4_42_108;
   wire n_4_42_109;
   wire n_4_42_110;
   wire n_4_42_111;
   wire n_4_42_112;
   wire n_4_42_113;
   wire n_4_42_114;
   wire n_4_42_115;
   wire n_4_42_116;
   wire n_4_42_117;
   wire n_4_42_118;
   wire n_4_42_119;
   wire n_4_42_120;
   wire n_4_42_121;
   wire n_4_42_122;
   wire n_4_42_123;
   wire n_4_42_124;
   wire n_4_42_125;
   wire n_4_42_126;
   wire n_4_42_127;
   wire n_4_42_128;
   wire n_4_42_129;
   wire n_4_42_130;
   wire n_4_42_131;
   wire n_4_42_132;
   wire n_4_42_133;
   wire n_4_42_134;
   wire n_4_42_135;
   wire n_4_42_136;
   wire n_4_42_137;
   wire n_4_42_138;
   wire n_4_42_139;
   wire n_4_42_140;
   wire n_4_42_141;
   wire n_4_42_142;
   wire n_4_42_143;
   wire n_4_42_144;
   wire n_5_41_0;
   wire n_5_41_1;
   wire n_5_41_2;
   wire n_5_41_3;
   wire n_5_41_4;
   wire n_5_41_5;
   wire n_5_41_6;
   wire n_5_41_7;
   wire n_5_41_8;
   wire n_5_41_9;
   wire n_5_41_10;
   wire n_5_41_11;
   wire n_5_41_12;
   wire n_5_41_13;
   wire n_5_41_14;
   wire n_5_41_15;
   wire n_5_41_16;
   wire n_5_41_17;
   wire n_5_41_18;
   wire n_5_41_19;
   wire n_5_41_20;
   wire n_5_41_21;
   wire n_5_41_22;
   wire n_5_41_23;
   wire n_5_41_24;
   wire n_5_41_25;
   wire n_5_41_26;
   wire n_5_41_27;
   wire n_5_41_28;
   wire n_5_41_29;
   wire n_5_41_30;
   wire n_5_41_31;
   wire n_5_41_32;
   wire n_5_41_33;
   wire n_5_41_34;
   wire n_5_41_35;
   wire n_5_41_36;
   wire n_5_41_37;
   wire n_5_41_38;
   wire n_5_41_39;
   wire n_5_41_40;
   wire n_5_41_41;
   wire n_5_41_42;
   wire n_5_41_43;
   wire n_5_41_44;
   wire n_5_41_45;
   wire n_5_41_46;
   wire n_5_41_47;
   wire n_5_41_48;
   wire n_5_41_49;
   wire n_5_41_50;
   wire n_5_41_51;
   wire n_5_41_52;
   wire n_5_41_53;
   wire n_5_41_54;
   wire n_5_41_55;
   wire n_5_41_56;
   wire n_5_41_57;
   wire n_5_41_58;
   wire n_5_41_59;
   wire n_5_41_60;
   wire n_5_41_61;
   wire n_5_41_62;
   wire n_5_41_63;
   wire n_5_41_64;
   wire n_5_41_65;
   wire n_5_41_66;
   wire n_5_41_67;
   wire n_5_41_68;
   wire n_5_41_69;
   wire n_5_41_70;
   wire n_5_41_71;
   wire n_5_41_72;
   wire n_5_41_73;
   wire n_5_41_74;
   wire n_5_41_75;
   wire n_5_41_76;
   wire n_5_41_77;
   wire n_5_41_78;
   wire n_5_41_79;
   wire n_5_41_80;
   wire n_5_41_81;
   wire n_5_41_82;
   wire n_5_41_83;
   wire n_5_41_84;
   wire n_5_41_85;
   wire n_5_41_86;
   wire n_5_41_87;
   wire n_5_41_88;
   wire n_5_41_89;
   wire n_5_41_90;
   wire n_5_41_91;
   wire n_5_41_92;
   wire n_5_41_93;
   wire n_5_41_94;
   wire n_5_41_95;
   wire n_5_41_96;
   wire n_5_41_97;
   wire n_5_41_98;
   wire n_5_41_99;
   wire n_5_41_100;
   wire n_5_41_101;
   wire n_5_41_102;
   wire n_5_41_103;
   wire n_5_41_104;
   wire n_5_41_105;
   wire n_5_41_106;
   wire n_5_41_107;
   wire n_5_41_108;
   wire n_5_41_109;
   wire n_5_41_110;
   wire n_5_41_111;
   wire n_5_41_112;
   wire n_5_41_113;
   wire n_5_41_114;
   wire n_5_41_115;
   wire n_5_41_116;
   wire n_5_41_117;
   wire n_5_41_118;
   wire n_5_41_119;
   wire n_5_41_120;
   wire n_5_41_121;
   wire n_5_41_122;
   wire n_5_41_123;
   wire n_5_41_124;
   wire n_5_41_125;
   wire n_5_41_126;
   wire n_5_41_127;
   wire n_5_41_128;
   wire n_5_41_129;
   wire n_5_41_130;
   wire n_5_41_131;
   wire n_5_41_132;
   wire n_5_41_133;
   wire n_5_41_134;
   wire n_5_41_135;
   wire n_5_41_136;
   wire n_5_41_137;
   wire n_5_41_138;
   wire n_5_41_139;
   wire n_5_41_140;
   wire n_5_41_141;
   wire n_5_41_142;
   wire n_5_41_143;
   wire n_5_41_144;
   wire n_6_40_0;
   wire n_6_40_1;
   wire n_6_40_2;
   wire n_6_40_3;
   wire n_6_40_4;
   wire n_6_40_5;
   wire n_6_40_6;
   wire n_6_40_7;
   wire n_6_40_8;
   wire n_6_40_9;
   wire n_6_40_10;
   wire n_6_40_11;
   wire n_6_40_12;
   wire n_6_40_13;
   wire n_6_40_14;
   wire n_6_40_15;
   wire n_6_40_16;
   wire n_6_40_17;
   wire n_6_40_18;
   wire n_6_40_19;
   wire n_6_40_20;
   wire n_6_40_21;
   wire n_6_40_22;
   wire n_6_40_23;
   wire n_6_40_24;
   wire n_6_40_25;
   wire n_6_40_26;
   wire n_6_40_27;
   wire n_6_40_28;
   wire n_6_40_29;
   wire n_6_40_30;
   wire n_6_40_31;
   wire n_6_40_32;
   wire n_6_40_33;
   wire n_6_40_34;
   wire n_6_40_35;
   wire n_6_40_36;
   wire n_6_40_37;
   wire n_6_40_38;
   wire n_6_40_39;
   wire n_6_40_40;
   wire n_6_40_41;
   wire n_6_40_42;
   wire n_6_40_43;
   wire n_6_40_44;
   wire n_6_40_45;
   wire n_6_40_46;
   wire n_6_40_47;
   wire n_6_40_48;
   wire n_6_40_49;
   wire n_6_40_50;
   wire n_6_40_51;
   wire n_6_40_52;
   wire n_6_40_53;
   wire n_6_40_54;
   wire n_6_40_55;
   wire n_6_40_56;
   wire n_6_40_57;
   wire n_6_40_58;
   wire n_6_40_59;
   wire n_6_40_60;
   wire n_6_40_61;
   wire n_6_40_62;
   wire n_6_40_63;
   wire n_6_40_64;
   wire n_6_40_65;
   wire n_6_40_66;
   wire n_6_40_67;
   wire n_6_40_68;
   wire n_6_40_69;
   wire n_6_40_70;
   wire n_6_40_71;
   wire n_6_40_72;
   wire n_6_40_73;
   wire n_6_40_74;
   wire n_6_40_75;
   wire n_6_40_76;
   wire n_6_40_77;
   wire n_6_40_78;
   wire n_6_40_79;
   wire n_6_40_80;
   wire n_6_40_81;
   wire n_6_40_82;
   wire n_6_40_83;
   wire n_6_40_84;
   wire n_6_40_85;
   wire n_6_40_86;
   wire n_6_40_87;
   wire n_6_40_88;
   wire n_6_40_89;
   wire n_6_40_90;
   wire n_6_40_91;
   wire n_6_40_92;
   wire n_6_40_93;
   wire n_6_40_94;
   wire n_6_40_95;
   wire n_6_40_96;
   wire n_6_40_97;
   wire n_6_40_98;
   wire n_6_40_99;
   wire n_6_40_100;
   wire n_6_40_101;
   wire n_6_40_102;
   wire n_6_40_103;
   wire n_6_40_104;
   wire n_6_40_105;
   wire n_6_40_106;
   wire n_6_40_107;
   wire n_6_40_108;
   wire n_6_40_109;
   wire n_6_40_110;
   wire n_6_40_111;
   wire n_6_40_112;
   wire n_6_40_113;
   wire n_6_40_114;
   wire n_6_40_115;
   wire n_6_40_116;
   wire n_6_40_117;
   wire n_6_40_118;
   wire n_6_40_119;
   wire n_6_40_120;
   wire n_6_40_121;
   wire n_6_40_122;
   wire n_6_40_123;
   wire n_6_40_124;
   wire n_6_40_125;
   wire n_6_40_126;
   wire n_6_40_127;
   wire n_6_40_128;
   wire n_6_40_129;
   wire n_6_40_130;
   wire n_6_40_131;
   wire n_6_40_132;
   wire n_6_40_133;
   wire n_6_40_134;
   wire n_6_40_135;
   wire n_6_40_136;
   wire n_6_40_137;
   wire n_6_40_138;
   wire n_6_40_139;
   wire n_6_40_140;
   wire n_6_40_141;
   wire n_6_40_142;
   wire n_6_40_143;
   wire n_6_40_144;
   wire n_7_39_0;
   wire n_7_39_1;
   wire n_7_39_2;
   wire n_7_39_3;
   wire n_7_39_4;
   wire n_7_39_5;
   wire n_7_39_6;
   wire n_7_39_7;
   wire n_7_39_8;
   wire n_7_39_9;
   wire n_7_39_10;
   wire n_7_39_11;
   wire n_7_39_12;
   wire n_7_39_13;
   wire n_7_39_14;
   wire n_7_39_15;
   wire n_7_39_16;
   wire n_7_39_17;
   wire n_7_39_18;
   wire n_7_39_19;
   wire n_7_39_20;
   wire n_7_39_21;
   wire n_7_39_22;
   wire n_7_39_23;
   wire n_7_39_24;
   wire n_7_39_25;
   wire n_7_39_26;
   wire n_7_39_27;
   wire n_7_39_28;
   wire n_7_39_29;
   wire n_7_39_30;
   wire n_7_39_31;
   wire n_7_39_32;
   wire n_7_39_33;
   wire n_7_39_34;
   wire n_7_39_35;
   wire n_7_39_36;
   wire n_7_39_37;
   wire n_7_39_38;
   wire n_7_39_39;
   wire n_7_39_40;
   wire n_7_39_41;
   wire n_7_39_42;
   wire n_7_39_43;
   wire n_7_39_44;
   wire n_7_39_45;
   wire n_7_39_46;
   wire n_7_39_47;
   wire n_7_39_48;
   wire n_7_39_49;
   wire n_7_39_50;
   wire n_7_39_51;
   wire n_7_39_52;
   wire n_7_39_53;
   wire n_7_39_54;
   wire n_7_39_55;
   wire n_7_39_56;
   wire n_7_39_57;
   wire n_7_39_58;
   wire n_7_39_59;
   wire n_7_39_60;
   wire n_7_39_61;
   wire n_7_39_62;
   wire n_7_39_63;
   wire n_7_39_64;
   wire n_7_39_65;
   wire n_7_39_66;
   wire n_7_39_67;
   wire n_7_39_68;
   wire n_7_39_69;
   wire n_7_39_70;
   wire n_7_39_71;
   wire n_7_39_72;
   wire n_7_39_73;
   wire n_7_39_74;
   wire n_7_39_75;
   wire n_7_39_76;
   wire n_7_39_77;
   wire n_7_39_78;
   wire n_7_39_79;
   wire n_7_39_80;
   wire n_7_39_81;
   wire n_7_39_82;
   wire n_7_39_83;
   wire n_7_39_84;
   wire n_7_39_85;
   wire n_7_39_86;
   wire n_7_39_87;
   wire n_7_39_88;
   wire n_7_39_89;
   wire n_7_39_90;
   wire n_7_39_91;
   wire n_7_39_92;
   wire n_7_39_93;
   wire n_7_39_94;
   wire n_7_39_95;
   wire n_7_39_96;
   wire n_7_39_97;
   wire n_7_39_98;
   wire n_7_39_99;
   wire n_7_39_100;
   wire n_7_39_101;
   wire n_7_39_102;
   wire n_7_39_103;
   wire n_7_39_104;
   wire n_7_39_105;
   wire n_7_39_106;
   wire n_7_39_107;
   wire n_7_39_108;
   wire n_7_39_109;
   wire n_7_39_110;
   wire n_7_39_111;
   wire n_7_39_112;
   wire n_7_39_113;
   wire n_7_39_114;
   wire n_7_39_115;
   wire n_7_39_116;
   wire n_7_39_117;
   wire n_7_39_118;
   wire n_7_39_119;
   wire n_7_39_120;
   wire n_7_39_121;
   wire n_7_39_122;
   wire n_7_39_123;
   wire n_7_39_124;
   wire n_7_39_125;
   wire n_7_39_126;
   wire n_7_39_127;
   wire n_7_39_128;
   wire n_7_39_129;
   wire n_7_39_130;
   wire n_7_39_131;
   wire n_7_39_132;
   wire n_7_39_133;
   wire n_7_39_134;
   wire n_7_39_135;
   wire n_7_39_136;
   wire n_7_39_137;
   wire n_7_39_138;
   wire n_7_39_139;
   wire n_7_39_140;
   wire n_7_39_141;
   wire n_7_39_142;
   wire n_7_39_143;
   wire n_7_39_144;
   wire n_8_37_0;
   wire n_8_37_1;
   wire n_8_37_2;
   wire n_8_37_3;
   wire n_8_37_4;
   wire n_8_37_5;
   wire n_8_37_6;
   wire n_8_37_7;
   wire n_8_37_8;
   wire n_8_37_9;
   wire n_8_37_10;
   wire n_8_37_11;
   wire n_8_37_12;
   wire n_8_37_13;
   wire n_8_37_14;
   wire n_8_37_15;
   wire n_8_37_16;
   wire n_8_37_17;
   wire n_8_37_18;
   wire n_8_37_19;
   wire n_8_37_20;
   wire n_8_37_21;
   wire n_8_37_22;
   wire n_8_37_23;
   wire n_8_37_24;
   wire n_8_37_25;
   wire n_8_37_26;
   wire n_8_37_27;
   wire n_8_37_28;
   wire n_8_37_29;
   wire n_8_37_30;
   wire n_8_37_31;
   wire n_8_37_32;
   wire n_8_37_33;
   wire n_8_37_34;
   wire n_8_37_35;
   wire n_8_37_36;
   wire n_8_37_37;
   wire n_8_37_38;
   wire n_8_37_39;
   wire n_8_37_40;
   wire n_8_37_41;
   wire n_8_37_42;
   wire n_8_37_43;
   wire n_8_37_44;
   wire n_8_37_45;
   wire n_8_37_46;
   wire n_8_37_47;
   wire n_8_37_48;
   wire n_8_37_49;
   wire n_8_37_50;
   wire n_8_37_51;
   wire n_8_37_52;
   wire n_8_37_53;
   wire n_8_37_54;
   wire n_8_37_55;
   wire n_8_37_56;
   wire n_8_37_57;
   wire n_8_37_58;
   wire n_8_37_59;
   wire n_8_37_60;
   wire n_8_37_61;
   wire n_8_37_62;
   wire n_8_37_63;
   wire n_8_37_64;
   wire n_8_37_65;
   wire n_8_37_66;
   wire n_8_37_67;
   wire n_8_37_68;
   wire n_8_37_69;
   wire n_8_37_70;
   wire n_8_37_71;
   wire n_8_37_72;
   wire n_8_37_73;
   wire n_8_37_74;
   wire n_8_37_75;
   wire n_8_37_76;
   wire n_8_37_77;
   wire n_8_37_78;
   wire n_8_37_79;
   wire n_8_37_80;
   wire n_8_37_81;
   wire n_8_37_82;
   wire n_8_37_83;
   wire n_8_37_84;
   wire n_8_37_85;
   wire n_8_37_86;
   wire n_8_37_87;
   wire n_8_37_88;
   wire n_8_37_89;
   wire n_8_37_90;
   wire n_8_37_91;
   wire n_8_37_92;
   wire n_8_37_93;
   wire n_8_37_94;
   wire n_8_37_95;
   wire n_8_37_96;
   wire n_8_37_97;
   wire n_8_37_98;
   wire n_8_37_99;
   wire n_8_37_100;
   wire n_8_37_101;
   wire n_8_37_102;
   wire n_8_37_103;
   wire n_8_37_104;
   wire n_8_37_105;
   wire n_8_37_106;
   wire n_8_37_107;
   wire n_8_37_108;
   wire n_8_37_109;
   wire n_8_37_110;
   wire n_8_37_111;
   wire n_8_37_112;
   wire n_8_37_113;
   wire n_8_37_114;
   wire n_8_37_115;
   wire n_8_37_116;
   wire n_8_37_117;
   wire n_8_37_118;
   wire n_8_37_119;
   wire n_8_37_120;
   wire n_8_37_121;
   wire n_8_37_122;
   wire n_8_37_123;
   wire n_8_37_124;
   wire n_8_37_125;
   wire n_8_37_126;
   wire n_8_37_127;
   wire n_8_37_128;
   wire n_8_37_129;
   wire n_8_37_130;
   wire n_8_37_131;
   wire n_8_37_132;
   wire n_8_37_133;
   wire n_8_37_134;
   wire n_8_37_135;
   wire n_8_37_136;
   wire n_8_37_137;
   wire n_8_37_138;
   wire n_8_37_139;
   wire n_8_37_140;
   wire n_8_37_141;
   wire n_8_37_142;
   wire n_8_37_143;
   wire n_8_37_144;
   wire n_9_36_0;
   wire n_9_36_1;
   wire n_9_36_2;
   wire n_9_36_3;
   wire n_9_36_4;
   wire n_9_36_5;
   wire n_9_36_6;
   wire n_9_36_7;
   wire n_9_36_8;
   wire n_9_36_9;
   wire n_9_36_10;
   wire n_9_36_11;
   wire n_9_36_12;
   wire n_9_36_13;
   wire n_9_36_14;
   wire n_9_36_15;
   wire n_9_36_16;
   wire n_9_36_17;
   wire n_9_36_18;
   wire n_9_36_19;
   wire n_9_36_20;
   wire n_9_36_21;
   wire n_9_36_22;
   wire n_9_36_23;
   wire n_9_36_24;
   wire n_9_36_25;
   wire n_9_36_26;
   wire n_9_36_27;
   wire n_9_36_28;
   wire n_9_36_29;
   wire n_9_36_30;
   wire n_9_36_31;
   wire n_9_36_32;
   wire n_9_36_33;
   wire n_9_36_34;
   wire n_9_36_35;
   wire n_9_36_36;
   wire n_9_36_37;
   wire n_9_36_38;
   wire n_9_36_39;
   wire n_9_36_40;
   wire n_9_36_41;
   wire n_9_36_42;
   wire n_9_36_43;
   wire n_9_36_44;
   wire n_9_36_45;
   wire n_9_36_46;
   wire n_9_36_47;
   wire n_9_36_48;
   wire n_9_36_49;
   wire n_9_36_50;
   wire n_9_36_51;
   wire n_9_36_52;
   wire n_9_36_53;
   wire n_9_36_54;
   wire n_9_36_55;
   wire n_9_36_56;
   wire n_9_36_57;
   wire n_9_36_58;
   wire n_9_36_59;
   wire n_9_36_60;
   wire n_9_36_61;
   wire n_9_36_62;
   wire n_9_36_63;
   wire n_9_36_64;
   wire n_9_36_65;
   wire n_9_36_66;
   wire n_9_36_67;
   wire n_9_36_68;
   wire n_9_36_69;
   wire n_9_36_70;
   wire n_9_36_71;
   wire n_9_36_72;
   wire n_9_36_73;
   wire n_9_36_74;
   wire n_9_36_75;
   wire n_9_36_76;
   wire n_9_36_77;
   wire n_9_36_78;
   wire n_9_36_79;
   wire n_9_36_80;
   wire n_9_36_81;
   wire n_9_36_82;
   wire n_9_36_83;
   wire n_9_36_84;
   wire n_9_36_85;
   wire n_9_36_86;
   wire n_9_36_87;
   wire n_9_36_88;
   wire n_9_36_89;
   wire n_9_36_90;
   wire n_9_36_91;
   wire n_9_36_92;
   wire n_9_36_93;
   wire n_9_36_94;
   wire n_9_36_95;
   wire n_9_36_96;
   wire n_9_36_97;
   wire n_9_36_98;
   wire n_9_36_99;
   wire n_9_36_100;
   wire n_9_36_101;
   wire n_9_36_102;
   wire n_9_36_103;
   wire n_9_36_104;
   wire n_9_36_105;
   wire n_9_36_106;
   wire n_9_36_107;
   wire n_9_36_108;
   wire n_9_36_109;
   wire n_9_36_110;
   wire n_9_36_111;
   wire n_9_36_112;
   wire n_9_36_113;
   wire n_9_36_114;
   wire n_9_36_115;
   wire n_9_36_116;
   wire n_9_36_117;
   wire n_9_36_118;
   wire n_9_36_119;
   wire n_9_36_120;
   wire n_9_36_121;
   wire n_9_36_122;
   wire n_9_36_123;
   wire n_9_36_124;
   wire n_9_36_125;
   wire n_9_36_126;
   wire n_9_36_127;
   wire n_9_36_128;
   wire n_9_36_129;
   wire n_9_36_130;
   wire n_9_36_131;
   wire n_9_36_132;
   wire n_9_36_133;
   wire n_9_36_134;
   wire n_9_36_135;
   wire n_9_36_136;
   wire n_9_36_137;
   wire n_9_36_138;
   wire n_9_36_139;
   wire n_9_36_140;
   wire n_9_36_141;
   wire n_9_36_142;
   wire n_9_36_143;
   wire n_9_36_144;
   wire n_10_35_0;
   wire n_10_35_1;
   wire n_10_35_2;
   wire n_10_35_3;
   wire n_10_35_4;
   wire n_10_35_5;
   wire n_10_35_6;
   wire n_10_35_7;
   wire n_10_35_8;
   wire n_10_35_9;
   wire n_10_35_10;
   wire n_10_35_11;
   wire n_10_35_12;
   wire n_10_35_13;
   wire n_10_35_14;
   wire n_10_35_15;
   wire n_10_35_16;
   wire n_10_35_17;
   wire n_10_35_18;
   wire n_10_35_19;
   wire n_10_35_20;
   wire n_10_35_21;
   wire n_10_35_22;
   wire n_10_35_23;
   wire n_10_35_24;
   wire n_10_35_25;
   wire n_10_35_26;
   wire n_10_35_27;
   wire n_10_35_28;
   wire n_10_35_29;
   wire n_10_35_30;
   wire n_10_35_31;
   wire n_10_35_32;
   wire n_10_35_33;
   wire n_10_35_34;
   wire n_10_35_35;
   wire n_10_35_36;
   wire n_10_35_37;
   wire n_10_35_38;
   wire n_10_35_39;
   wire n_10_35_40;
   wire n_10_35_41;
   wire n_10_35_42;
   wire n_10_35_43;
   wire n_10_35_44;
   wire n_10_35_45;
   wire n_10_35_46;
   wire n_10_35_47;
   wire n_10_35_48;
   wire n_10_35_49;
   wire n_10_35_50;
   wire n_10_35_51;
   wire n_10_35_52;
   wire n_10_35_53;
   wire n_10_35_54;
   wire n_10_35_55;
   wire n_10_35_56;
   wire n_10_35_57;
   wire n_10_35_58;
   wire n_10_35_59;
   wire n_10_35_60;
   wire n_10_35_61;
   wire n_10_35_62;
   wire n_10_35_63;
   wire n_10_35_64;
   wire n_10_35_65;
   wire n_10_35_66;
   wire n_10_35_67;
   wire n_10_35_68;
   wire n_10_35_69;
   wire n_10_35_70;
   wire n_10_35_71;
   wire n_10_35_72;
   wire n_10_35_73;
   wire n_10_35_74;
   wire n_10_35_75;
   wire n_10_35_76;
   wire n_10_35_77;
   wire n_10_35_78;
   wire n_10_35_79;
   wire n_10_35_80;
   wire n_10_35_81;
   wire n_10_35_82;
   wire n_10_35_83;
   wire n_10_35_84;
   wire n_10_35_85;
   wire n_10_35_86;
   wire n_10_35_87;
   wire n_10_35_88;
   wire n_10_35_89;
   wire n_10_35_90;
   wire n_10_35_91;
   wire n_10_35_92;
   wire n_10_35_93;
   wire n_10_35_94;
   wire n_10_35_95;
   wire n_10_35_96;
   wire n_10_35_97;
   wire n_10_35_98;
   wire n_10_35_99;
   wire n_10_35_100;
   wire n_10_35_101;
   wire n_10_35_102;
   wire n_10_35_103;
   wire n_10_35_104;
   wire n_10_35_105;
   wire n_10_35_106;
   wire n_10_35_107;
   wire n_10_35_108;
   wire n_10_35_109;
   wire n_10_35_110;
   wire n_10_35_111;
   wire n_10_35_112;
   wire n_10_35_113;
   wire n_10_35_114;
   wire n_10_35_115;
   wire n_10_35_116;
   wire n_10_35_117;
   wire n_10_35_118;
   wire n_10_35_119;
   wire n_10_35_120;
   wire n_10_35_121;
   wire n_10_35_122;
   wire n_10_35_123;
   wire n_10_35_124;
   wire n_10_35_125;
   wire n_10_35_126;
   wire n_10_35_127;
   wire n_10_35_128;
   wire n_10_35_129;
   wire n_10_35_130;
   wire n_10_35_131;
   wire n_10_35_132;
   wire n_10_35_133;
   wire n_10_35_134;
   wire n_10_35_135;
   wire n_10_35_136;
   wire n_10_35_137;
   wire n_10_35_138;
   wire n_10_35_139;
   wire n_10_35_140;
   wire n_10_35_141;
   wire n_10_35_142;
   wire n_10_35_143;
   wire n_10_35_144;
   wire n_11_33_0;
   wire n_11_33_1;
   wire n_11_33_2;
   wire n_11_33_3;
   wire n_11_33_4;
   wire n_11_33_5;
   wire n_11_33_6;
   wire n_11_33_7;
   wire n_11_33_8;
   wire n_11_33_9;
   wire n_11_33_10;
   wire n_11_33_11;
   wire n_11_33_12;
   wire n_11_33_13;
   wire n_11_33_14;
   wire n_11_33_15;
   wire n_11_33_16;
   wire n_11_33_17;
   wire n_11_33_18;
   wire n_11_33_19;
   wire n_11_33_20;
   wire n_11_33_21;
   wire n_11_33_22;
   wire n_11_33_23;
   wire n_11_33_24;
   wire n_11_33_25;
   wire n_11_33_26;
   wire n_11_33_27;
   wire n_11_33_28;
   wire n_11_33_29;
   wire n_11_33_30;
   wire n_11_33_31;
   wire n_11_33_32;
   wire n_11_33_33;
   wire n_11_33_34;
   wire n_11_33_35;
   wire n_11_33_36;
   wire n_11_33_37;
   wire n_11_33_38;
   wire n_11_33_39;
   wire n_11_33_40;
   wire n_11_33_41;
   wire n_11_33_42;
   wire n_11_33_43;
   wire n_11_33_44;
   wire n_11_33_45;
   wire n_11_33_46;
   wire n_11_33_47;
   wire n_11_33_48;
   wire n_11_33_49;
   wire n_11_33_50;
   wire n_11_33_51;
   wire n_11_33_52;
   wire n_11_33_53;
   wire n_11_33_54;
   wire n_11_33_55;
   wire n_11_33_56;
   wire n_11_33_57;
   wire n_11_33_58;
   wire n_11_33_59;
   wire n_11_33_60;
   wire n_11_33_61;
   wire n_11_33_62;
   wire n_11_33_63;
   wire n_11_33_64;
   wire n_11_33_65;
   wire n_11_33_66;
   wire n_11_33_67;
   wire n_11_33_68;
   wire n_11_33_69;
   wire n_11_33_70;
   wire n_11_33_71;
   wire n_11_33_72;
   wire n_11_33_73;
   wire n_11_33_74;
   wire n_11_33_75;
   wire n_11_33_76;
   wire n_11_33_77;
   wire n_11_33_78;
   wire n_11_33_79;
   wire n_11_33_80;
   wire n_11_33_81;
   wire n_11_33_82;
   wire n_11_33_83;
   wire n_11_33_84;
   wire n_11_33_85;
   wire n_11_33_86;
   wire n_11_33_87;
   wire n_11_33_88;
   wire n_11_33_89;
   wire n_11_33_90;
   wire n_11_33_91;
   wire n_11_33_92;
   wire n_11_33_93;
   wire n_11_33_94;
   wire n_11_33_95;
   wire n_11_33_96;
   wire n_11_33_97;
   wire n_11_33_98;
   wire n_11_33_99;
   wire n_11_33_100;
   wire n_11_33_101;
   wire n_11_33_102;
   wire n_11_33_103;
   wire n_11_33_104;
   wire n_11_33_105;
   wire n_11_33_106;
   wire n_11_33_107;
   wire n_11_33_108;
   wire n_11_33_109;
   wire n_11_33_110;
   wire n_11_33_111;
   wire n_11_33_112;
   wire n_11_33_113;
   wire n_11_33_114;
   wire n_11_33_115;
   wire n_11_33_116;
   wire n_11_33_117;
   wire n_11_33_118;
   wire n_11_33_119;
   wire n_11_33_120;
   wire n_11_33_121;
   wire n_11_33_122;
   wire n_11_33_123;
   wire n_11_33_124;
   wire n_11_33_125;
   wire n_11_33_126;
   wire n_11_33_127;
   wire n_11_33_128;
   wire n_11_33_129;
   wire n_11_33_130;
   wire n_11_33_131;
   wire n_11_33_132;
   wire n_11_33_133;
   wire n_11_33_134;
   wire n_11_33_135;
   wire n_11_33_136;
   wire n_11_33_137;
   wire n_11_33_138;
   wire n_11_33_139;
   wire n_11_33_140;
   wire n_11_33_141;
   wire n_11_33_142;
   wire n_11_33_143;
   wire n_11_33_144;
   wire n_12_32_0;
   wire n_12_32_1;
   wire n_12_32_2;
   wire n_12_32_3;
   wire n_12_32_4;
   wire n_12_32_5;
   wire n_12_32_6;
   wire n_12_32_7;
   wire n_12_32_8;
   wire n_12_32_9;
   wire n_12_32_10;
   wire n_12_32_11;
   wire n_12_32_12;
   wire n_12_32_13;
   wire n_12_32_14;
   wire n_12_32_15;
   wire n_12_32_16;
   wire n_12_32_17;
   wire n_12_32_18;
   wire n_12_32_19;
   wire n_12_32_20;
   wire n_12_32_21;
   wire n_12_32_22;
   wire n_12_32_23;
   wire n_12_32_24;
   wire n_12_32_25;
   wire n_12_32_26;
   wire n_12_32_27;
   wire n_12_32_28;
   wire n_12_32_29;
   wire n_12_32_30;
   wire n_12_32_31;
   wire n_12_32_32;
   wire n_12_32_33;
   wire n_12_32_34;
   wire n_12_32_35;
   wire n_12_32_36;
   wire n_12_32_37;
   wire n_12_32_38;
   wire n_12_32_39;
   wire n_12_32_40;
   wire n_12_32_41;
   wire n_12_32_42;
   wire n_12_32_43;
   wire n_12_32_44;
   wire n_12_32_45;
   wire n_12_32_46;
   wire n_12_32_47;
   wire n_12_32_48;
   wire n_12_32_49;
   wire n_12_32_50;
   wire n_12_32_51;
   wire n_12_32_52;
   wire n_12_32_53;
   wire n_12_32_54;
   wire n_12_32_55;
   wire n_12_32_56;
   wire n_12_32_57;
   wire n_12_32_58;
   wire n_12_32_59;
   wire n_12_32_60;
   wire n_12_32_61;
   wire n_12_32_62;
   wire n_12_32_63;
   wire n_12_32_64;
   wire n_12_32_65;
   wire n_12_32_66;
   wire n_12_32_67;
   wire n_12_32_68;
   wire n_12_32_69;
   wire n_12_32_70;
   wire n_12_32_71;
   wire n_12_32_72;
   wire n_12_32_73;
   wire n_12_32_74;
   wire n_12_32_75;
   wire n_12_32_76;
   wire n_12_32_77;
   wire n_12_32_78;
   wire n_12_32_79;
   wire n_12_32_80;
   wire n_12_32_81;
   wire n_12_32_82;
   wire n_12_32_83;
   wire n_12_32_84;
   wire n_12_32_85;
   wire n_12_32_86;
   wire n_12_32_87;
   wire n_12_32_88;
   wire n_12_32_89;
   wire n_12_32_90;
   wire n_12_32_91;
   wire n_12_32_92;
   wire n_12_32_93;
   wire n_12_32_94;
   wire n_12_32_95;
   wire n_12_32_96;
   wire n_12_32_97;
   wire n_12_32_98;
   wire n_12_32_99;
   wire n_12_32_100;
   wire n_12_32_101;
   wire n_12_32_102;
   wire n_12_32_103;
   wire n_12_32_104;
   wire n_12_32_105;
   wire n_12_32_106;
   wire n_12_32_107;
   wire n_12_32_108;
   wire n_12_32_109;
   wire n_12_32_110;
   wire n_12_32_111;
   wire n_12_32_112;
   wire n_12_32_113;
   wire n_12_32_114;
   wire n_12_32_115;
   wire n_12_32_116;
   wire n_12_32_117;
   wire n_12_32_118;
   wire n_12_32_119;
   wire n_12_32_120;
   wire n_12_32_121;
   wire n_12_32_122;
   wire n_12_32_123;
   wire n_12_32_124;
   wire n_12_32_125;
   wire n_12_32_126;
   wire n_12_32_127;
   wire n_12_32_128;
   wire n_12_32_129;
   wire n_12_32_130;
   wire n_12_32_131;
   wire n_12_32_132;
   wire n_12_32_133;
   wire n_12_32_134;
   wire n_12_32_135;
   wire n_12_32_136;
   wire n_12_32_137;
   wire n_12_32_138;
   wire n_12_32_139;
   wire n_12_32_140;
   wire n_12_32_141;
   wire n_12_32_142;
   wire n_12_32_143;
   wire n_12_32_144;
   wire n_13_31_0;
   wire n_13_31_1;
   wire n_13_31_2;
   wire n_13_31_3;
   wire n_13_31_4;
   wire n_13_31_5;
   wire n_13_31_6;
   wire n_13_31_7;
   wire n_13_31_8;
   wire n_13_31_9;
   wire n_13_31_10;
   wire n_13_31_11;
   wire n_13_31_12;
   wire n_13_31_13;
   wire n_13_31_14;
   wire n_13_31_15;
   wire n_13_31_16;
   wire n_13_31_17;
   wire n_13_31_18;
   wire n_13_31_19;
   wire n_13_31_20;
   wire n_13_31_21;
   wire n_13_31_22;
   wire n_13_31_23;
   wire n_13_31_24;
   wire n_13_31_25;
   wire n_13_31_26;
   wire n_13_31_27;
   wire n_13_31_28;
   wire n_13_31_29;
   wire n_13_31_30;
   wire n_13_31_31;
   wire n_13_31_32;
   wire n_13_31_33;
   wire n_13_31_34;
   wire n_13_31_35;
   wire n_13_31_36;
   wire n_13_31_37;
   wire n_13_31_38;
   wire n_13_31_39;
   wire n_13_31_40;
   wire n_13_31_41;
   wire n_13_31_42;
   wire n_13_31_43;
   wire n_13_31_44;
   wire n_13_31_45;
   wire n_13_31_46;
   wire n_13_31_47;
   wire n_13_31_48;
   wire n_13_31_49;
   wire n_13_31_50;
   wire n_13_31_51;
   wire n_13_31_52;
   wire n_13_31_53;
   wire n_13_31_54;
   wire n_13_31_55;
   wire n_13_31_56;
   wire n_13_31_57;
   wire n_13_31_58;
   wire n_13_31_59;
   wire n_13_31_60;
   wire n_13_31_61;
   wire n_13_31_62;
   wire n_13_31_63;
   wire n_13_31_64;
   wire n_13_31_65;
   wire n_13_31_66;
   wire n_13_31_67;
   wire n_13_31_68;
   wire n_13_31_69;
   wire n_13_31_70;
   wire n_13_31_71;
   wire n_13_31_72;
   wire n_13_31_73;
   wire n_13_31_74;
   wire n_13_31_75;
   wire n_13_31_76;
   wire n_13_31_77;
   wire n_13_31_78;
   wire n_13_31_79;
   wire n_13_31_80;
   wire n_13_31_81;
   wire n_13_31_82;
   wire n_13_31_83;
   wire n_13_31_84;
   wire n_13_31_85;
   wire n_13_31_86;
   wire n_13_31_87;
   wire n_13_31_88;
   wire n_13_31_89;
   wire n_13_31_90;
   wire n_13_31_91;
   wire n_13_31_92;
   wire n_13_31_93;
   wire n_13_31_94;
   wire n_13_31_95;
   wire n_13_31_96;
   wire n_13_31_97;
   wire n_13_31_98;
   wire n_13_31_99;
   wire n_13_31_100;
   wire n_13_31_101;
   wire n_13_31_102;
   wire n_13_31_103;
   wire n_13_31_104;
   wire n_13_31_105;
   wire n_13_31_106;
   wire n_13_31_107;
   wire n_13_31_108;
   wire n_13_31_109;
   wire n_13_31_110;
   wire n_13_31_111;
   wire n_13_31_112;
   wire n_13_31_113;
   wire n_13_31_114;
   wire n_13_31_115;
   wire n_13_31_116;
   wire n_13_31_117;
   wire n_13_31_118;
   wire n_13_31_119;
   wire n_13_31_120;
   wire n_13_31_121;
   wire n_13_31_122;
   wire n_13_31_123;
   wire n_13_31_124;
   wire n_13_31_125;
   wire n_13_31_126;
   wire n_13_31_127;
   wire n_13_31_128;
   wire n_13_31_129;
   wire n_13_31_130;
   wire n_13_31_131;
   wire n_13_31_132;
   wire n_13_31_133;
   wire n_13_31_134;
   wire n_13_31_135;
   wire n_13_31_136;
   wire n_13_31_137;
   wire n_13_31_138;
   wire n_13_31_139;
   wire n_13_31_140;
   wire n_13_31_141;
   wire n_13_31_142;
   wire n_13_31_143;
   wire n_13_31_144;
   wire n_14_30_0;
   wire n_14_30_1;
   wire n_14_30_2;
   wire n_14_30_3;
   wire n_14_30_4;
   wire n_14_30_5;
   wire n_14_30_6;
   wire n_14_30_7;
   wire n_14_30_8;
   wire n_14_30_9;
   wire n_14_30_10;
   wire n_14_30_11;
   wire n_14_30_12;
   wire n_14_30_13;
   wire n_14_30_14;
   wire n_14_30_15;
   wire n_14_30_16;
   wire n_14_30_17;
   wire n_14_30_18;
   wire n_14_30_19;
   wire n_14_30_20;
   wire n_14_30_21;
   wire n_14_30_22;
   wire n_14_30_23;
   wire n_14_30_24;
   wire n_14_30_25;
   wire n_14_30_26;
   wire n_14_30_27;
   wire n_14_30_28;
   wire n_14_30_29;
   wire n_14_30_30;
   wire n_14_30_31;
   wire n_14_30_32;
   wire n_14_30_33;
   wire n_14_30_34;
   wire n_14_30_35;
   wire n_14_30_36;
   wire n_14_30_37;
   wire n_14_30_38;
   wire n_14_30_39;
   wire n_14_30_40;
   wire n_14_30_41;
   wire n_14_30_42;
   wire n_14_30_43;
   wire n_14_30_44;
   wire n_14_30_45;
   wire n_14_30_46;
   wire n_14_30_47;
   wire n_14_30_48;
   wire n_14_30_49;
   wire n_14_30_50;
   wire n_14_30_51;
   wire n_14_30_52;
   wire n_14_30_53;
   wire n_14_30_54;
   wire n_14_30_55;
   wire n_14_30_56;
   wire n_14_30_57;
   wire n_14_30_58;
   wire n_14_30_59;
   wire n_14_30_60;
   wire n_14_30_61;
   wire n_14_30_62;
   wire n_14_30_63;
   wire n_14_30_64;
   wire n_14_30_65;
   wire n_14_30_66;
   wire n_14_30_67;
   wire n_14_30_68;
   wire n_14_30_69;
   wire n_14_30_70;
   wire n_14_30_71;
   wire n_14_30_72;
   wire n_14_30_73;
   wire n_14_30_74;
   wire n_14_30_75;
   wire n_14_30_76;
   wire n_14_30_77;
   wire n_14_30_78;
   wire n_14_30_79;
   wire n_14_30_80;
   wire n_14_30_81;
   wire n_14_30_82;
   wire n_14_30_83;
   wire n_14_30_84;
   wire n_14_30_85;
   wire n_14_30_86;
   wire n_14_30_87;
   wire n_14_30_88;
   wire n_14_30_89;
   wire n_14_30_90;
   wire n_14_30_91;
   wire n_14_30_92;
   wire n_14_30_93;
   wire n_14_30_94;
   wire n_14_30_95;
   wire n_14_30_96;
   wire n_14_30_97;
   wire n_14_30_98;
   wire n_14_30_99;
   wire n_14_30_100;
   wire n_14_30_101;
   wire n_14_30_102;
   wire n_14_30_103;
   wire n_14_30_104;
   wire n_14_30_105;
   wire n_14_30_106;
   wire n_14_30_107;
   wire n_14_30_108;
   wire n_14_30_109;
   wire n_14_30_110;
   wire n_14_30_111;
   wire n_14_30_112;
   wire n_14_30_113;
   wire n_14_30_114;
   wire n_14_30_115;
   wire n_14_30_116;
   wire n_14_30_117;
   wire n_14_30_118;
   wire n_14_30_119;
   wire n_14_30_120;
   wire n_14_30_121;
   wire n_14_30_122;
   wire n_14_30_123;
   wire n_14_30_124;
   wire n_14_30_125;
   wire n_14_30_126;
   wire n_14_30_127;
   wire n_14_30_128;
   wire n_14_30_129;
   wire n_14_30_130;
   wire n_14_30_131;
   wire n_14_30_132;
   wire n_14_30_133;
   wire n_14_30_134;
   wire n_14_30_135;
   wire n_14_30_136;
   wire n_14_30_137;
   wire n_14_30_138;
   wire n_14_30_139;
   wire n_14_30_140;
   wire n_14_30_141;
   wire n_14_30_142;
   wire n_14_30_143;
   wire n_14_30_144;
   wire n_15_29_0;
   wire n_15_29_1;
   wire n_15_29_2;
   wire n_15_29_3;
   wire n_15_29_4;
   wire n_15_29_5;
   wire n_15_29_6;
   wire n_15_29_7;
   wire n_15_29_8;
   wire n_15_29_9;
   wire n_15_29_10;
   wire n_15_29_11;
   wire n_15_29_12;
   wire n_15_29_13;
   wire n_15_29_14;
   wire n_15_29_15;
   wire n_15_29_16;
   wire n_15_29_17;
   wire n_15_29_18;
   wire n_15_29_19;
   wire n_15_29_20;
   wire n_15_29_21;
   wire n_15_29_22;
   wire n_15_29_23;
   wire n_15_29_24;
   wire n_15_29_25;
   wire n_15_29_26;
   wire n_15_29_27;
   wire n_15_29_28;
   wire n_15_29_29;
   wire n_15_29_30;
   wire n_15_29_31;
   wire n_15_29_32;
   wire n_15_29_33;
   wire n_15_29_34;
   wire n_15_29_35;
   wire n_15_29_36;
   wire n_15_29_37;
   wire n_15_29_38;
   wire n_15_29_39;
   wire n_15_29_40;
   wire n_15_29_41;
   wire n_15_29_42;
   wire n_15_29_43;
   wire n_15_29_44;
   wire n_15_29_45;
   wire n_15_29_46;
   wire n_15_29_47;
   wire n_15_29_48;
   wire n_15_29_49;
   wire n_15_29_50;
   wire n_15_29_51;
   wire n_15_29_52;
   wire n_15_29_53;
   wire n_15_29_54;
   wire n_15_29_55;
   wire n_15_29_56;
   wire n_15_29_57;
   wire n_15_29_58;
   wire n_15_29_59;
   wire n_15_29_60;
   wire n_15_29_61;
   wire n_15_29_62;
   wire n_15_29_63;
   wire n_15_29_64;
   wire n_15_29_65;
   wire n_15_29_66;
   wire n_15_29_67;
   wire n_15_29_68;
   wire n_15_29_69;
   wire n_15_29_70;
   wire n_15_29_71;
   wire n_15_29_72;
   wire n_15_29_73;
   wire n_15_29_74;
   wire n_15_29_75;
   wire n_15_29_76;
   wire n_15_29_77;
   wire n_15_29_78;
   wire n_15_29_79;
   wire n_15_29_80;
   wire n_15_29_81;
   wire n_15_29_82;
   wire n_15_29_83;
   wire n_15_29_84;
   wire n_15_29_85;
   wire n_15_29_86;
   wire n_15_29_87;
   wire n_15_29_88;
   wire n_15_29_89;
   wire n_15_29_90;
   wire n_15_29_91;
   wire n_15_29_92;
   wire n_15_29_93;
   wire n_15_29_94;
   wire n_15_29_95;
   wire n_15_29_96;
   wire n_15_29_97;
   wire n_15_29_98;
   wire n_15_29_99;
   wire n_15_29_100;
   wire n_15_29_101;
   wire n_15_29_102;
   wire n_15_29_103;
   wire n_15_29_104;
   wire n_15_29_105;
   wire n_15_29_106;
   wire n_15_29_107;
   wire n_15_29_108;
   wire n_15_29_109;
   wire n_15_29_110;
   wire n_15_29_111;
   wire n_15_29_112;
   wire n_15_29_113;
   wire n_15_29_114;
   wire n_15_29_115;
   wire n_15_29_116;
   wire n_15_29_117;
   wire n_15_29_118;
   wire n_15_29_119;
   wire n_15_29_120;
   wire n_15_29_121;
   wire n_15_29_122;
   wire n_15_29_123;
   wire n_15_29_124;
   wire n_15_29_125;
   wire n_15_29_126;
   wire n_15_29_127;
   wire n_15_29_128;
   wire n_15_29_129;
   wire n_15_29_130;
   wire n_15_29_131;
   wire n_15_29_132;
   wire n_15_29_133;
   wire n_15_29_134;
   wire n_15_29_135;
   wire n_15_29_136;
   wire n_15_29_137;
   wire n_15_29_138;
   wire n_15_29_139;
   wire n_15_29_140;
   wire n_15_29_141;
   wire n_15_29_142;
   wire n_15_29_143;
   wire n_15_29_144;
   wire n_16_28_0;
   wire n_16_28_1;
   wire n_16_28_2;
   wire n_16_28_3;
   wire n_16_28_4;
   wire n_16_28_5;
   wire n_16_28_6;
   wire n_16_28_7;
   wire n_16_28_8;
   wire n_16_28_9;
   wire n_16_28_10;
   wire n_16_28_11;
   wire n_16_28_12;
   wire n_16_28_13;
   wire n_16_28_14;
   wire n_16_28_15;
   wire n_16_28_16;
   wire n_16_28_17;
   wire n_16_28_18;
   wire n_16_28_19;
   wire n_16_28_20;
   wire n_16_28_21;
   wire n_16_28_22;
   wire n_16_28_23;
   wire n_16_28_24;
   wire n_16_28_25;
   wire n_16_28_26;
   wire n_16_28_27;
   wire n_16_28_28;
   wire n_16_28_29;
   wire n_16_28_30;
   wire n_16_28_31;
   wire n_16_28_32;
   wire n_16_28_33;
   wire n_16_28_34;
   wire n_16_28_35;
   wire n_16_28_36;
   wire n_16_28_37;
   wire n_16_28_38;
   wire n_16_28_39;
   wire n_16_28_40;
   wire n_16_28_41;
   wire n_16_28_42;
   wire n_16_28_43;
   wire n_16_28_44;
   wire n_16_28_45;
   wire n_16_28_46;
   wire n_16_28_47;
   wire n_16_28_48;
   wire n_16_28_49;
   wire n_16_28_50;
   wire n_16_28_51;
   wire n_16_28_52;
   wire n_16_28_53;
   wire n_16_28_54;
   wire n_16_28_55;
   wire n_16_28_56;
   wire n_16_28_57;
   wire n_16_28_58;
   wire n_16_28_59;
   wire n_16_28_60;
   wire n_16_28_61;
   wire n_16_28_62;
   wire n_16_28_63;
   wire n_16_28_64;
   wire n_16_28_65;
   wire n_16_28_66;
   wire n_16_28_67;
   wire n_16_28_68;
   wire n_16_28_69;
   wire n_16_28_70;
   wire n_16_28_71;
   wire n_16_28_72;
   wire n_16_28_73;
   wire n_16_28_74;
   wire n_16_28_75;
   wire n_16_28_76;
   wire n_16_28_77;
   wire n_16_28_78;
   wire n_16_28_79;
   wire n_16_28_80;
   wire n_16_28_81;
   wire n_16_28_82;
   wire n_16_28_83;
   wire n_16_28_84;
   wire n_16_28_85;
   wire n_16_28_86;
   wire n_16_28_87;
   wire n_16_28_88;
   wire n_16_28_89;
   wire n_16_28_90;
   wire n_16_28_91;
   wire n_16_28_92;
   wire n_16_28_93;
   wire n_16_28_94;
   wire n_16_28_95;
   wire n_16_28_96;
   wire n_16_28_97;
   wire n_16_28_98;
   wire n_16_28_99;
   wire n_16_28_100;
   wire n_16_28_101;
   wire n_16_28_102;
   wire n_16_28_103;
   wire n_16_28_104;
   wire n_16_28_105;
   wire n_16_28_106;
   wire n_16_28_107;
   wire n_16_28_108;
   wire n_16_28_109;
   wire n_16_28_110;
   wire n_16_28_111;
   wire n_16_28_112;
   wire n_16_28_113;
   wire n_16_28_114;
   wire n_16_28_115;
   wire n_16_28_116;
   wire n_16_28_117;
   wire n_16_28_118;
   wire n_16_28_119;
   wire n_16_28_120;
   wire n_16_28_121;
   wire n_16_28_122;
   wire n_16_28_123;
   wire n_16_28_124;
   wire n_16_28_125;
   wire n_16_28_126;
   wire n_16_28_127;
   wire n_16_28_128;
   wire n_16_28_129;
   wire n_16_28_130;
   wire n_16_28_131;
   wire n_16_28_132;
   wire n_16_28_133;
   wire n_16_28_134;
   wire n_16_28_135;
   wire n_16_28_136;
   wire n_16_28_137;
   wire n_16_28_138;
   wire n_16_28_139;
   wire n_16_28_140;
   wire n_16_28_141;
   wire n_16_28_142;
   wire n_16_28_143;
   wire n_16_28_144;
   wire n_17_34_0;
   wire n_17_34_1;
   wire n_17_34_2;
   wire n_17_34_3;
   wire n_17_34_4;
   wire n_17_34_5;
   wire n_17_34_6;
   wire n_17_34_7;
   wire n_17_34_8;
   wire n_17_34_9;
   wire n_17_34_10;
   wire n_17_34_11;
   wire n_17_34_12;
   wire n_17_34_13;
   wire n_17_34_14;
   wire n_17_34_15;
   wire n_17_34_16;
   wire n_17_34_17;
   wire n_17_34_18;
   wire n_17_34_19;
   wire n_17_34_20;
   wire n_17_34_21;
   wire n_17_34_22;
   wire n_17_34_23;
   wire n_17_34_24;
   wire n_17_34_25;
   wire n_17_34_26;
   wire n_17_34_27;
   wire n_17_34_28;
   wire n_17_34_29;
   wire n_17_34_30;
   wire n_17_34_31;
   wire n_17_34_32;
   wire n_17_34_33;
   wire n_17_34_34;
   wire n_17_34_35;
   wire n_17_34_36;
   wire n_17_34_37;
   wire n_17_34_38;
   wire n_17_34_39;
   wire n_17_34_40;
   wire n_17_34_41;
   wire n_17_34_42;
   wire n_17_34_43;
   wire n_17_34_44;
   wire n_17_34_45;
   wire n_17_34_46;
   wire n_17_34_47;
   wire n_17_34_48;
   wire n_17_34_49;
   wire n_17_34_50;
   wire n_17_34_51;
   wire n_17_34_52;
   wire n_17_34_53;
   wire n_17_34_54;
   wire n_17_34_55;
   wire n_17_34_56;
   wire n_17_34_57;
   wire n_17_34_58;
   wire n_17_34_59;
   wire n_17_34_60;
   wire n_17_34_61;
   wire n_17_34_62;
   wire n_17_34_63;
   wire n_17_34_64;
   wire n_17_34_65;
   wire n_17_34_66;
   wire n_17_34_67;
   wire n_17_34_68;
   wire n_17_34_69;
   wire n_17_34_70;
   wire n_17_34_71;
   wire n_17_34_72;
   wire n_17_34_73;
   wire n_17_34_74;
   wire n_17_34_75;
   wire n_17_34_76;
   wire n_17_34_77;
   wire n_17_34_78;
   wire n_17_34_79;
   wire n_17_34_80;
   wire n_17_34_81;
   wire n_17_34_82;
   wire n_17_34_83;
   wire n_17_34_84;
   wire n_17_34_85;
   wire n_17_34_86;
   wire n_17_34_87;
   wire n_17_34_88;
   wire n_17_34_89;
   wire n_17_34_90;
   wire n_17_34_91;
   wire n_17_34_92;
   wire n_17_34_93;
   wire n_17_34_94;
   wire n_17_34_95;
   wire n_17_34_96;
   wire n_17_34_97;
   wire n_17_34_98;
   wire n_17_34_99;
   wire n_17_34_100;
   wire n_17_34_101;
   wire n_17_34_102;
   wire n_17_34_103;
   wire n_17_34_104;
   wire n_17_34_105;
   wire n_17_34_106;
   wire n_17_34_107;
   wire n_17_34_108;
   wire n_17_34_109;
   wire n_17_34_110;
   wire n_17_34_111;
   wire n_17_34_112;
   wire n_17_34_113;
   wire n_17_34_114;
   wire n_17_34_115;
   wire n_17_34_116;
   wire n_17_34_117;
   wire n_17_34_118;
   wire n_17_34_119;
   wire n_17_34_120;
   wire n_17_34_121;
   wire n_17_34_122;
   wire n_17_34_123;
   wire n_17_34_124;
   wire n_17_34_125;
   wire n_17_34_126;
   wire n_17_34_127;
   wire n_17_34_128;
   wire n_17_34_129;
   wire n_17_34_130;
   wire n_17_34_131;
   wire n_17_34_132;
   wire n_17_34_133;
   wire n_17_34_134;
   wire n_17_34_135;
   wire n_17_34_136;
   wire n_17_34_137;
   wire n_17_34_138;
   wire n_17_34_139;
   wire n_17_34_140;
   wire n_17_34_141;
   wire n_17_34_142;
   wire n_17_34_143;
   wire n_17_34_144;
   wire n_27_27_0;
   wire n_27_27_1;
   wire n_27_27_2;
   wire n_27_27_3;
   wire n_27_27_4;
   wire n_27_27_5;
   wire n_27_27_6;
   wire n_27_27_7;
   wire n_27_27_8;
   wire n_27_27_9;
   wire n_27_27_10;
   wire n_27_27_11;
   wire n_27_27_12;
   wire n_27_27_13;
   wire n_27_27_14;
   wire n_27_27_15;
   wire n_27_27_16;
   wire n_27_27_17;
   wire n_27_27_18;
   wire n_27_27_19;
   wire n_27_27_20;
   wire n_27_27_21;
   wire n_27_27_22;
   wire n_27_27_23;
   wire n_27_27_24;
   wire n_27_27_25;
   wire n_27_27_26;
   wire n_27_27_27;
   wire n_27_27_28;
   wire n_27_27_29;
   wire n_27_27_30;
   wire n_27_27_31;
   wire n_27_27_32;
   wire n_27_27_33;
   wire n_27_27_34;
   wire n_27_27_35;
   wire n_27_27_36;
   wire n_27_27_37;
   wire n_27_27_38;
   wire n_27_27_39;
   wire n_27_27_40;
   wire n_27_27_41;
   wire n_27_27_42;
   wire n_27_27_43;
   wire n_27_27_44;
   wire n_27_27_45;
   wire n_27_27_46;
   wire n_27_27_47;
   wire n_27_27_48;
   wire n_27_27_49;
   wire n_27_27_50;
   wire n_27_27_51;
   wire n_27_27_52;
   wire n_27_27_53;
   wire n_27_27_54;
   wire n_27_27_55;
   wire n_27_27_56;
   wire n_27_27_57;
   wire n_27_27_58;
   wire n_27_27_59;
   wire n_27_27_60;
   wire n_27_27_61;
   wire n_27_27_62;
   wire n_27_27_63;
   wire n_27_27_64;
   wire n_27_27_65;
   wire n_27_27_66;
   wire n_27_27_67;
   wire n_27_27_68;
   wire n_27_27_69;
   wire n_27_27_70;
   wire n_27_27_71;
   wire n_27_27_72;
   wire n_27_27_73;
   wire n_27_27_74;
   wire n_27_27_75;
   wire n_27_27_76;
   wire n_27_27_77;
   wire n_27_27_78;
   wire n_27_27_79;
   wire n_27_27_80;
   wire n_27_27_81;
   wire n_27_27_82;
   wire n_27_27_83;
   wire n_27_27_84;
   wire n_27_27_85;
   wire n_27_27_86;
   wire n_27_27_87;
   wire n_27_27_88;
   wire n_27_27_89;
   wire n_27_27_90;
   wire n_27_27_91;
   wire n_27_27_92;
   wire n_27_27_93;
   wire n_27_27_94;
   wire n_27_27_95;
   wire n_27_27_96;
   wire n_27_27_97;
   wire n_27_27_98;
   wire n_27_27_99;
   wire n_27_27_100;
   wire n_27_27_101;
   wire n_27_27_102;
   wire n_27_27_103;
   wire n_27_27_104;
   wire n_27_27_105;
   wire n_27_27_106;
   wire n_27_27_107;
   wire n_27_27_108;
   wire n_27_27_109;
   wire n_27_27_110;
   wire n_27_27_111;
   wire n_27_27_112;
   wire n_27_27_113;
   wire n_27_27_114;
   wire n_27_27_115;
   wire n_27_27_116;
   wire n_27_27_117;
   wire n_27_27_118;
   wire n_27_27_119;
   wire n_27_27_120;
   wire n_27_27_121;
   wire n_27_27_122;
   wire n_27_27_123;
   wire n_27_27_124;
   wire n_27_27_125;
   wire n_27_27_126;
   wire n_27_27_127;
   wire n_27_27_128;
   wire n_27_27_129;
   wire n_27_27_130;
   wire n_27_27_131;
   wire n_27_27_132;
   wire n_27_27_133;
   wire n_27_27_134;
   wire n_27_27_135;
   wire n_27_27_136;
   wire n_27_27_137;
   wire n_27_27_138;
   wire n_27_27_139;
   wire n_27_27_140;
   wire n_27_27_141;
   wire n_27_27_142;
   wire n_27_27_143;
   wire n_27_27_144;
   wire n_26_26_0;
   wire n_26_26_1;
   wire n_26_26_2;
   wire n_26_26_3;
   wire n_26_26_4;
   wire n_26_26_5;
   wire n_26_26_6;
   wire n_26_26_7;
   wire n_26_26_8;
   wire n_26_26_9;
   wire n_26_26_10;
   wire n_26_26_11;
   wire n_26_26_12;
   wire n_26_26_13;
   wire n_26_26_14;
   wire n_26_26_15;
   wire n_26_26_16;
   wire n_26_26_17;
   wire n_26_26_18;
   wire n_26_26_19;
   wire n_26_26_20;
   wire n_26_26_21;
   wire n_26_26_22;
   wire n_26_26_23;
   wire n_26_26_24;
   wire n_26_26_25;
   wire n_26_26_26;
   wire n_26_26_27;
   wire n_26_26_28;
   wire n_26_26_29;
   wire n_26_26_30;
   wire n_26_26_31;
   wire n_26_26_32;
   wire n_26_26_33;
   wire n_26_26_34;
   wire n_26_26_35;
   wire n_26_26_36;
   wire n_26_26_37;
   wire n_26_26_38;
   wire n_26_26_39;
   wire n_26_26_40;
   wire n_26_26_41;
   wire n_26_26_42;
   wire n_26_26_43;
   wire n_26_26_44;
   wire n_26_26_45;
   wire n_26_26_46;
   wire n_26_26_47;
   wire n_26_26_48;
   wire n_26_26_49;
   wire n_26_26_50;
   wire n_26_26_51;
   wire n_26_26_52;
   wire n_26_26_53;
   wire n_26_26_54;
   wire n_26_26_55;
   wire n_26_26_56;
   wire n_26_26_57;
   wire n_26_26_58;
   wire n_26_26_59;
   wire n_26_26_60;
   wire n_26_26_61;
   wire n_26_26_62;
   wire n_26_26_63;
   wire n_26_26_64;
   wire n_26_26_65;
   wire n_26_26_66;
   wire n_26_26_67;
   wire n_26_26_68;
   wire n_26_26_69;
   wire n_26_26_70;
   wire n_26_26_71;
   wire n_26_26_72;
   wire n_26_26_73;
   wire n_26_26_74;
   wire n_26_26_75;
   wire n_26_26_76;
   wire n_26_26_77;
   wire n_26_26_78;
   wire n_26_26_79;
   wire n_26_26_80;
   wire n_26_26_81;
   wire n_26_26_82;
   wire n_26_26_83;
   wire n_26_26_84;
   wire n_26_26_85;
   wire n_26_26_86;
   wire n_26_26_87;
   wire n_26_26_88;
   wire n_26_26_89;
   wire n_26_26_90;
   wire n_26_26_91;
   wire n_26_26_92;
   wire n_26_26_93;
   wire n_26_26_94;
   wire n_26_26_95;
   wire n_26_26_96;
   wire n_26_26_97;
   wire n_26_26_98;
   wire n_26_26_99;
   wire n_26_26_100;
   wire n_26_26_101;
   wire n_26_26_102;
   wire n_26_26_103;
   wire n_26_26_104;
   wire n_26_26_105;
   wire n_26_26_106;
   wire n_26_26_107;
   wire n_26_26_108;
   wire n_26_26_109;
   wire n_26_26_110;
   wire n_26_26_111;
   wire n_26_26_112;
   wire n_26_26_113;
   wire n_26_26_114;
   wire n_26_26_115;
   wire n_26_26_116;
   wire n_26_26_117;
   wire n_26_26_118;
   wire n_26_26_119;
   wire n_26_26_120;
   wire n_26_26_121;
   wire n_26_26_122;
   wire n_26_26_123;
   wire n_26_26_124;
   wire n_26_26_125;
   wire n_26_26_126;
   wire n_26_26_127;
   wire n_26_26_128;
   wire n_26_26_129;
   wire n_26_26_130;
   wire n_26_26_131;
   wire n_26_26_132;
   wire n_26_26_133;
   wire n_26_26_134;
   wire n_26_26_135;
   wire n_26_26_136;
   wire n_26_26_137;
   wire n_26_26_138;
   wire n_26_26_139;
   wire n_26_26_140;
   wire n_26_26_141;
   wire n_26_26_142;
   wire n_26_26_143;
   wire n_26_26_144;
   wire n_25_25_0;
   wire n_25_25_1;
   wire n_25_25_2;
   wire n_25_25_3;
   wire n_25_25_4;
   wire n_25_25_5;
   wire n_25_25_6;
   wire n_25_25_7;
   wire n_25_25_8;
   wire n_25_25_9;
   wire n_25_25_10;
   wire n_25_25_11;
   wire n_25_25_12;
   wire n_25_25_13;
   wire n_25_25_14;
   wire n_25_25_15;
   wire n_25_25_16;
   wire n_25_25_17;
   wire n_25_25_18;
   wire n_25_25_19;
   wire n_25_25_20;
   wire n_25_25_21;
   wire n_25_25_22;
   wire n_25_25_23;
   wire n_25_25_24;
   wire n_25_25_25;
   wire n_25_25_26;
   wire n_25_25_27;
   wire n_25_25_28;
   wire n_25_25_29;
   wire n_25_25_30;
   wire n_25_25_31;
   wire n_25_25_32;
   wire n_25_25_33;
   wire n_25_25_34;
   wire n_25_25_35;
   wire n_25_25_36;
   wire n_25_25_37;
   wire n_25_25_38;
   wire n_25_25_39;
   wire n_25_25_40;
   wire n_25_25_41;
   wire n_25_25_42;
   wire n_25_25_43;
   wire n_25_25_44;
   wire n_25_25_45;
   wire n_25_25_46;
   wire n_25_25_47;
   wire n_25_25_48;
   wire n_25_25_49;
   wire n_25_25_50;
   wire n_25_25_51;
   wire n_25_25_52;
   wire n_25_25_53;
   wire n_25_25_54;
   wire n_25_25_55;
   wire n_25_25_56;
   wire n_25_25_57;
   wire n_25_25_58;
   wire n_25_25_59;
   wire n_25_25_60;
   wire n_25_25_61;
   wire n_25_25_62;
   wire n_25_25_63;
   wire n_25_25_64;
   wire n_25_25_65;
   wire n_25_25_66;
   wire n_25_25_67;
   wire n_25_25_68;
   wire n_25_25_69;
   wire n_25_25_70;
   wire n_25_25_71;
   wire n_25_25_72;
   wire n_25_25_73;
   wire n_25_25_74;
   wire n_25_25_75;
   wire n_25_25_76;
   wire n_25_25_77;
   wire n_25_25_78;
   wire n_25_25_79;
   wire n_25_25_80;
   wire n_25_25_81;
   wire n_25_25_82;
   wire n_25_25_83;
   wire n_25_25_84;
   wire n_25_25_85;
   wire n_25_25_86;
   wire n_25_25_87;
   wire n_25_25_88;
   wire n_25_25_89;
   wire n_25_25_90;
   wire n_25_25_91;
   wire n_25_25_92;
   wire n_25_25_93;
   wire n_25_25_94;
   wire n_25_25_95;
   wire n_25_25_96;
   wire n_25_25_97;
   wire n_25_25_98;
   wire n_25_25_99;
   wire n_25_25_100;
   wire n_25_25_101;
   wire n_25_25_102;
   wire n_25_25_103;
   wire n_25_25_104;
   wire n_25_25_105;
   wire n_25_25_106;
   wire n_25_25_107;
   wire n_25_25_108;
   wire n_25_25_109;
   wire n_25_25_110;
   wire n_25_25_111;
   wire n_25_25_112;
   wire n_25_25_113;
   wire n_25_25_114;
   wire n_25_25_115;
   wire n_25_25_116;
   wire n_25_25_117;
   wire n_25_25_118;
   wire n_25_25_119;
   wire n_25_25_120;
   wire n_25_25_121;
   wire n_25_25_122;
   wire n_25_25_123;
   wire n_25_25_124;
   wire n_25_25_125;
   wire n_25_25_126;
   wire n_25_25_127;
   wire n_25_25_128;
   wire n_25_25_129;
   wire n_25_25_130;
   wire n_25_25_131;
   wire n_25_25_132;
   wire n_25_25_133;
   wire n_25_25_134;
   wire n_25_25_135;
   wire n_25_25_136;
   wire n_25_25_137;
   wire n_25_25_138;
   wire n_25_25_139;
   wire n_25_25_140;
   wire n_25_25_141;
   wire n_25_25_142;
   wire n_25_25_143;
   wire n_25_25_144;
   wire n_28_38_0;
   wire n_28_38_1;
   wire n_28_38_2;
   wire n_28_38_3;
   wire n_28_38_4;
   wire n_28_38_5;
   wire n_28_38_6;
   wire n_28_38_7;
   wire n_28_38_8;
   wire n_28_38_9;
   wire n_28_38_10;
   wire n_28_38_11;
   wire n_28_38_12;
   wire n_28_38_13;
   wire n_28_38_14;
   wire n_28_38_15;
   wire n_28_38_16;
   wire n_28_38_17;
   wire n_28_38_18;
   wire n_28_38_19;
   wire n_28_38_20;
   wire n_28_38_21;
   wire n_28_38_22;
   wire n_28_38_23;
   wire n_28_38_24;
   wire n_28_38_25;
   wire n_28_38_26;
   wire n_28_38_27;
   wire n_28_38_28;
   wire n_28_38_29;
   wire n_28_38_30;
   wire n_28_38_31;
   wire n_28_38_32;
   wire n_28_38_33;
   wire n_28_38_34;
   wire n_28_38_35;
   wire n_28_38_36;
   wire n_28_38_37;
   wire n_28_38_38;
   wire n_28_38_39;
   wire n_28_38_40;
   wire n_28_38_41;
   wire n_28_38_42;
   wire n_28_38_43;
   wire n_28_38_44;
   wire n_28_38_45;
   wire n_28_38_46;
   wire n_28_38_47;
   wire n_28_38_48;
   wire n_28_38_49;
   wire n_28_38_50;
   wire n_28_38_51;
   wire n_28_38_52;
   wire n_28_38_53;
   wire n_28_38_54;
   wire n_28_38_55;
   wire n_28_38_56;
   wire n_28_38_57;
   wire n_28_38_58;
   wire n_28_38_59;
   wire n_28_38_60;
   wire n_28_38_61;
   wire n_28_38_62;
   wire n_28_38_63;
   wire n_28_38_64;
   wire n_28_38_65;
   wire n_28_38_66;
   wire n_28_38_67;
   wire n_28_38_68;
   wire n_28_38_69;
   wire n_28_38_70;
   wire n_28_38_71;
   wire n_28_38_72;
   wire n_28_38_73;
   wire n_28_38_74;
   wire n_28_38_75;
   wire n_28_38_76;
   wire n_28_38_77;
   wire n_28_38_78;
   wire n_28_38_79;
   wire n_28_38_80;
   wire n_28_38_81;
   wire n_28_38_82;
   wire n_28_38_83;
   wire n_28_38_84;
   wire n_28_38_85;
   wire n_28_38_86;
   wire n_28_38_87;
   wire n_28_38_88;
   wire n_28_38_89;
   wire n_28_38_90;
   wire n_28_38_91;
   wire n_28_38_92;
   wire n_28_38_93;
   wire n_28_38_94;
   wire n_28_38_95;
   wire n_28_38_96;
   wire n_28_38_97;
   wire n_28_38_98;
   wire n_28_38_99;
   wire n_28_38_100;
   wire n_28_38_101;
   wire n_28_38_102;
   wire n_28_38_103;
   wire n_28_38_104;
   wire n_28_38_105;
   wire n_28_38_106;
   wire n_28_38_107;
   wire n_28_38_108;
   wire n_28_38_109;
   wire n_28_38_110;
   wire n_28_38_111;
   wire n_28_38_112;
   wire n_28_38_113;
   wire n_28_38_114;
   wire n_28_38_115;
   wire n_28_38_116;
   wire n_28_38_117;
   wire n_28_38_118;
   wire n_28_38_119;
   wire n_28_38_120;
   wire n_28_38_121;
   wire n_28_38_122;
   wire n_28_38_123;
   wire n_28_38_124;
   wire n_28_38_125;
   wire n_28_38_126;
   wire n_28_38_127;
   wire n_28_38_128;
   wire n_28_38_129;
   wire n_28_38_130;
   wire n_28_38_131;
   wire n_28_38_132;
   wire n_28_38_133;
   wire n_28_38_134;
   wire n_28_38_135;
   wire n_28_38_136;
   wire n_28_38_137;
   wire n_28_38_138;
   wire n_28_38_139;
   wire n_28_38_140;
   wire n_28_38_141;
   wire n_28_38_142;
   wire n_28_38_143;
   wire n_28_38_144;
   wire n_24_24_0;
   wire n_24_24_1;
   wire n_24_24_2;
   wire n_24_24_3;
   wire n_24_24_4;
   wire n_24_24_5;
   wire n_24_24_6;
   wire n_24_24_7;
   wire n_24_24_8;
   wire n_24_24_9;
   wire n_24_24_10;
   wire n_24_24_11;
   wire n_24_24_12;
   wire n_24_24_13;
   wire n_24_24_14;
   wire n_24_24_15;
   wire n_24_24_16;
   wire n_24_24_17;
   wire n_24_24_18;
   wire n_24_24_19;
   wire n_24_24_20;
   wire n_24_24_21;
   wire n_24_24_22;
   wire n_24_24_23;
   wire n_24_24_24;
   wire n_24_24_25;
   wire n_24_24_26;
   wire n_24_24_27;
   wire n_24_24_28;
   wire n_24_24_29;
   wire n_24_24_30;
   wire n_24_24_31;
   wire n_24_24_32;
   wire n_24_24_33;
   wire n_24_24_34;
   wire n_24_24_35;
   wire n_24_24_36;
   wire n_24_24_37;
   wire n_24_24_38;
   wire n_24_24_39;
   wire n_24_24_40;
   wire n_24_24_41;
   wire n_24_24_42;
   wire n_24_24_43;
   wire n_24_24_44;
   wire n_24_24_45;
   wire n_24_24_46;
   wire n_24_24_47;
   wire n_24_24_48;
   wire n_24_24_49;
   wire n_24_24_50;
   wire n_24_24_51;
   wire n_24_24_52;
   wire n_24_24_53;
   wire n_24_24_54;
   wire n_24_24_55;
   wire n_24_24_56;
   wire n_24_24_57;
   wire n_24_24_58;
   wire n_24_24_59;
   wire n_24_24_60;
   wire n_24_24_61;
   wire n_24_24_62;
   wire n_24_24_63;
   wire n_24_24_64;
   wire n_24_24_65;
   wire n_24_24_66;
   wire n_24_24_67;
   wire n_24_24_68;
   wire n_24_24_69;
   wire n_24_24_70;
   wire n_24_24_71;
   wire n_24_24_72;
   wire n_24_24_73;
   wire n_24_24_74;
   wire n_24_24_75;
   wire n_24_24_76;
   wire n_24_24_77;
   wire n_24_24_78;
   wire n_24_24_79;
   wire n_24_24_80;
   wire n_24_24_81;
   wire n_24_24_82;
   wire n_24_24_83;
   wire n_24_24_84;
   wire n_24_24_85;
   wire n_24_24_86;
   wire n_24_24_87;
   wire n_24_24_88;
   wire n_24_24_89;
   wire n_24_24_90;
   wire n_24_24_91;
   wire n_24_24_92;
   wire n_24_24_93;
   wire n_24_24_94;
   wire n_24_24_95;
   wire n_24_24_96;
   wire n_24_24_97;
   wire n_24_24_98;
   wire n_24_24_99;
   wire n_24_24_100;
   wire n_24_24_101;
   wire n_24_24_102;
   wire n_24_24_103;
   wire n_24_24_104;
   wire n_24_24_105;
   wire n_24_24_106;
   wire n_24_24_107;
   wire n_24_24_108;
   wire n_24_24_109;
   wire n_24_24_110;
   wire n_24_24_111;
   wire n_24_24_112;
   wire n_24_24_113;
   wire n_24_24_114;
   wire n_24_24_115;
   wire n_24_24_116;
   wire n_24_24_117;
   wire n_24_24_118;
   wire n_24_24_119;
   wire n_24_24_120;
   wire n_24_24_121;
   wire n_24_24_122;
   wire n_24_24_123;
   wire n_24_24_124;
   wire n_24_24_125;
   wire n_24_24_126;
   wire n_24_24_127;
   wire n_24_24_128;
   wire n_24_24_129;
   wire n_24_24_130;
   wire n_24_24_131;
   wire n_24_24_132;
   wire n_24_24_133;
   wire n_24_24_134;
   wire n_24_24_135;
   wire n_24_24_136;
   wire n_24_24_137;
   wire n_24_24_138;
   wire n_24_24_139;
   wire n_24_24_140;
   wire n_24_24_141;
   wire n_24_24_142;
   wire n_24_24_143;
   wire n_24_24_144;
   wire n_23_23_0;
   wire n_23_23_1;
   wire n_23_23_2;
   wire n_23_23_3;
   wire n_23_23_4;
   wire n_23_23_5;
   wire n_23_23_6;
   wire n_23_23_7;
   wire n_23_23_8;
   wire n_23_23_9;
   wire n_23_23_10;
   wire n_23_23_11;
   wire n_23_23_12;
   wire n_23_23_13;
   wire n_23_23_14;
   wire n_23_23_15;
   wire n_23_23_16;
   wire n_23_23_17;
   wire n_23_23_18;
   wire n_23_23_19;
   wire n_23_23_20;
   wire n_23_23_21;
   wire n_23_23_22;
   wire n_23_23_23;
   wire n_23_23_24;
   wire n_23_23_25;
   wire n_23_23_26;
   wire n_23_23_27;
   wire n_23_23_28;
   wire n_23_23_29;
   wire n_23_23_30;
   wire n_23_23_31;
   wire n_23_23_32;
   wire n_23_23_33;
   wire n_23_23_34;
   wire n_23_23_35;
   wire n_23_23_36;
   wire n_23_23_37;
   wire n_23_23_38;
   wire n_23_23_39;
   wire n_23_23_40;
   wire n_23_23_41;
   wire n_23_23_42;
   wire n_23_23_43;
   wire n_23_23_44;
   wire n_23_23_45;
   wire n_23_23_46;
   wire n_23_23_47;
   wire n_23_23_48;
   wire n_23_23_49;
   wire n_23_23_50;
   wire n_23_23_51;
   wire n_23_23_52;
   wire n_23_23_53;
   wire n_23_23_54;
   wire n_23_23_55;
   wire n_23_23_56;
   wire n_23_23_57;
   wire n_23_23_58;
   wire n_23_23_59;
   wire n_23_23_60;
   wire n_23_23_61;
   wire n_23_23_62;
   wire n_23_23_63;
   wire n_23_23_64;
   wire n_23_23_65;
   wire n_23_23_66;
   wire n_23_23_67;
   wire n_23_23_68;
   wire n_23_23_69;
   wire n_23_23_70;
   wire n_23_23_71;
   wire n_23_23_72;
   wire n_23_23_73;
   wire n_23_23_74;
   wire n_23_23_75;
   wire n_23_23_76;
   wire n_23_23_77;
   wire n_23_23_78;
   wire n_23_23_79;
   wire n_23_23_80;
   wire n_23_23_81;
   wire n_23_23_82;
   wire n_23_23_83;
   wire n_23_23_84;
   wire n_23_23_85;
   wire n_23_23_86;
   wire n_23_23_87;
   wire n_23_23_88;
   wire n_23_23_89;
   wire n_23_23_90;
   wire n_23_23_91;
   wire n_23_23_92;
   wire n_23_23_93;
   wire n_23_23_94;
   wire n_23_23_95;
   wire n_23_23_96;
   wire n_23_23_97;
   wire n_23_23_98;
   wire n_23_23_99;
   wire n_23_23_100;
   wire n_23_23_101;
   wire n_23_23_102;
   wire n_23_23_103;
   wire n_23_23_104;
   wire n_23_23_105;
   wire n_23_23_106;
   wire n_23_23_107;
   wire n_23_23_108;
   wire n_23_23_109;
   wire n_23_23_110;
   wire n_23_23_111;
   wire n_23_23_112;
   wire n_23_23_113;
   wire n_23_23_114;
   wire n_23_23_115;
   wire n_23_23_116;
   wire n_23_23_117;
   wire n_23_23_118;
   wire n_23_23_119;
   wire n_23_23_120;
   wire n_23_23_121;
   wire n_23_23_122;
   wire n_23_23_123;
   wire n_23_23_124;
   wire n_23_23_125;
   wire n_23_23_126;
   wire n_23_23_127;
   wire n_23_23_128;
   wire n_23_23_129;
   wire n_23_23_130;
   wire n_23_23_131;
   wire n_23_23_132;
   wire n_23_23_133;
   wire n_23_23_134;
   wire n_23_23_135;
   wire n_23_23_136;
   wire n_23_23_137;
   wire n_23_23_138;
   wire n_23_23_139;
   wire n_23_23_140;
   wire n_23_23_141;
   wire n_23_23_142;
   wire n_23_23_143;
   wire n_23_23_144;
   wire n_22_22_0;
   wire n_22_22_1;
   wire n_22_22_2;
   wire n_22_22_3;
   wire n_22_22_4;
   wire n_22_22_5;
   wire n_22_22_6;
   wire n_22_22_7;
   wire n_22_22_8;
   wire n_22_22_9;
   wire n_22_22_10;
   wire n_22_22_11;
   wire n_22_22_12;
   wire n_22_22_13;
   wire n_22_22_14;
   wire n_22_22_15;
   wire n_22_22_16;
   wire n_22_22_17;
   wire n_22_22_18;
   wire n_22_22_19;
   wire n_22_22_20;
   wire n_22_22_21;
   wire n_22_22_22;
   wire n_22_22_23;
   wire n_22_22_24;
   wire n_22_22_25;
   wire n_22_22_26;
   wire n_22_22_27;
   wire n_22_22_28;
   wire n_22_22_29;
   wire n_22_22_30;
   wire n_22_22_31;
   wire n_22_22_32;
   wire n_22_22_33;
   wire n_22_22_34;
   wire n_22_22_35;
   wire n_22_22_36;
   wire n_22_22_37;
   wire n_22_22_38;
   wire n_22_22_39;
   wire n_22_22_40;
   wire n_22_22_41;
   wire n_22_22_42;
   wire n_22_22_43;
   wire n_22_22_44;
   wire n_22_22_45;
   wire n_22_22_46;
   wire n_22_22_47;
   wire n_22_22_48;
   wire n_22_22_49;
   wire n_22_22_50;
   wire n_22_22_51;
   wire n_22_22_52;
   wire n_22_22_53;
   wire n_22_22_54;
   wire n_22_22_55;
   wire n_22_22_56;
   wire n_22_22_57;
   wire n_22_22_58;
   wire n_22_22_59;
   wire n_22_22_60;
   wire n_22_22_61;
   wire n_22_22_62;
   wire n_22_22_63;
   wire n_22_22_64;
   wire n_22_22_65;
   wire n_22_22_66;
   wire n_22_22_67;
   wire n_22_22_68;
   wire n_22_22_69;
   wire n_22_22_70;
   wire n_22_22_71;
   wire n_22_22_72;
   wire n_22_22_73;
   wire n_22_22_74;
   wire n_22_22_75;
   wire n_22_22_76;
   wire n_22_22_77;
   wire n_22_22_78;
   wire n_22_22_79;
   wire n_22_22_80;
   wire n_22_22_81;
   wire n_22_22_82;
   wire n_22_22_83;
   wire n_22_22_84;
   wire n_22_22_85;
   wire n_22_22_86;
   wire n_22_22_87;
   wire n_22_22_88;
   wire n_22_22_89;
   wire n_22_22_90;
   wire n_22_22_91;
   wire n_22_22_92;
   wire n_22_22_93;
   wire n_22_22_94;
   wire n_22_22_95;
   wire n_22_22_96;
   wire n_22_22_97;
   wire n_22_22_98;
   wire n_22_22_99;
   wire n_22_22_100;
   wire n_22_22_101;
   wire n_22_22_102;
   wire n_22_22_103;
   wire n_22_22_104;
   wire n_22_22_105;
   wire n_22_22_106;
   wire n_22_22_107;
   wire n_22_22_108;
   wire n_22_22_109;
   wire n_22_22_110;
   wire n_22_22_111;
   wire n_22_22_112;
   wire n_22_22_113;
   wire n_22_22_114;
   wire n_22_22_115;
   wire n_22_22_116;
   wire n_22_22_117;
   wire n_22_22_118;
   wire n_22_22_119;
   wire n_22_22_120;
   wire n_22_22_121;
   wire n_22_22_122;
   wire n_22_22_123;
   wire n_22_22_124;
   wire n_22_22_125;
   wire n_22_22_126;
   wire n_22_22_127;
   wire n_22_22_128;
   wire n_22_22_129;
   wire n_22_22_130;
   wire n_22_22_131;
   wire n_22_22_132;
   wire n_22_22_133;
   wire n_22_22_134;
   wire n_22_22_135;
   wire n_22_22_136;
   wire n_22_22_137;
   wire n_22_22_138;
   wire n_22_22_139;
   wire n_22_22_140;
   wire n_22_22_141;
   wire n_22_22_142;
   wire n_22_22_143;
   wire n_22_22_144;
   wire n_21_21_0;
   wire n_21_21_1;
   wire n_21_21_2;
   wire n_21_21_3;
   wire n_21_21_4;
   wire n_21_21_5;
   wire n_21_21_6;
   wire n_21_21_7;
   wire n_21_21_8;
   wire n_21_21_9;
   wire n_21_21_10;
   wire n_21_21_11;
   wire n_21_21_12;
   wire n_21_21_13;
   wire n_21_21_14;
   wire n_21_21_15;
   wire n_21_21_16;
   wire n_21_21_17;
   wire n_21_21_18;
   wire n_21_21_19;
   wire n_21_21_20;
   wire n_21_21_21;
   wire n_21_21_22;
   wire n_21_21_23;
   wire n_21_21_24;
   wire n_21_21_25;
   wire n_21_21_26;
   wire n_21_21_27;
   wire n_21_21_28;
   wire n_21_21_29;
   wire n_21_21_30;
   wire n_21_21_31;
   wire n_21_21_32;
   wire n_21_21_33;
   wire n_21_21_34;
   wire n_21_21_35;
   wire n_21_21_36;
   wire n_21_21_37;
   wire n_21_21_38;
   wire n_21_21_39;
   wire n_21_21_40;
   wire n_21_21_41;
   wire n_21_21_42;
   wire n_21_21_43;
   wire n_21_21_44;
   wire n_21_21_45;
   wire n_21_21_46;
   wire n_21_21_47;
   wire n_21_21_48;
   wire n_21_21_49;
   wire n_21_21_50;
   wire n_21_21_51;
   wire n_21_21_52;
   wire n_21_21_53;
   wire n_21_21_54;
   wire n_21_21_55;
   wire n_21_21_56;
   wire n_21_21_57;
   wire n_21_21_58;
   wire n_21_21_59;
   wire n_21_21_60;
   wire n_21_21_61;
   wire n_21_21_62;
   wire n_21_21_63;
   wire n_21_21_64;
   wire n_21_21_65;
   wire n_21_21_66;
   wire n_21_21_67;
   wire n_21_21_68;
   wire n_21_21_69;
   wire n_21_21_70;
   wire n_21_21_71;
   wire n_21_21_72;
   wire n_21_21_73;
   wire n_21_21_74;
   wire n_21_21_75;
   wire n_21_21_76;
   wire n_21_21_77;
   wire n_21_21_78;
   wire n_21_21_79;
   wire n_21_21_80;
   wire n_21_21_81;
   wire n_21_21_82;
   wire n_21_21_83;
   wire n_21_21_84;
   wire n_21_21_85;
   wire n_21_21_86;
   wire n_21_21_87;
   wire n_21_21_88;
   wire n_21_21_89;
   wire n_21_21_90;
   wire n_21_21_91;
   wire n_21_21_92;
   wire n_21_21_93;
   wire n_21_21_94;
   wire n_21_21_95;
   wire n_21_21_96;
   wire n_21_21_97;
   wire n_21_21_98;
   wire n_21_21_99;
   wire n_21_21_100;
   wire n_21_21_101;
   wire n_21_21_102;
   wire n_21_21_103;
   wire n_21_21_104;
   wire n_21_21_105;
   wire n_21_21_106;
   wire n_21_21_107;
   wire n_21_21_108;
   wire n_21_21_109;
   wire n_21_21_110;
   wire n_21_21_111;
   wire n_21_21_112;
   wire n_21_21_113;
   wire n_21_21_114;
   wire n_21_21_115;
   wire n_21_21_116;
   wire n_21_21_117;
   wire n_21_21_118;
   wire n_21_21_119;
   wire n_21_21_120;
   wire n_21_21_121;
   wire n_21_21_122;
   wire n_21_21_123;
   wire n_21_21_124;
   wire n_21_21_125;
   wire n_21_21_126;
   wire n_21_21_127;
   wire n_21_21_128;
   wire n_21_21_129;
   wire n_21_21_130;
   wire n_21_21_131;
   wire n_21_21_132;
   wire n_21_21_133;
   wire n_21_21_134;
   wire n_21_21_135;
   wire n_21_21_136;
   wire n_21_21_137;
   wire n_21_21_138;
   wire n_21_21_139;
   wire n_21_21_140;
   wire n_21_21_141;
   wire n_21_21_142;
   wire n_21_21_143;
   wire n_21_21_144;
   wire n_19_0_0;
   wire n_19_0_1;
   wire n_19_0_2;
   wire n_19_0_3;
   wire n_19_0_4;
   wire n_19_0_5;
   wire n_19_0_6;
   wire n_19_0_7;
   wire n_19_0_8;
   wire n_19_0_9;
   wire n_19_0_10;
   wire n_19_0_11;
   wire n_19_0_12;
   wire n_19_0_13;
   wire n_19_0_14;
   wire n_19_0_15;
   wire n_19_0_16;
   wire n_19_0_17;
   wire n_19_0_18;
   wire n_19_0_19;
   wire n_19_0_20;
   wire n_19_0_21;
   wire n_19_0_22;
   wire n_19_0_23;
   wire n_19_0_24;
   wire n_19_0_25;
   wire n_19_0_26;
   wire n_19_0_27;
   wire n_19_0_28;
   wire n_19_0_29;
   wire n_19_0_30;
   wire n_19_0_31;
   wire n_19_0_32;
   wire n_19_0_33;
   wire n_19_0_34;
   wire n_19_0_35;
   wire n_19_0_36;
   wire n_19_0_37;
   wire n_19_0_38;
   wire n_19_0_39;
   wire n_19_0_40;
   wire n_19_0_41;
   wire n_19_0_42;
   wire n_19_0_43;
   wire n_19_0_44;
   wire n_19_0_45;
   wire n_19_0_46;
   wire n_19_0_47;
   wire n_19_0_48;
   wire n_19_0_49;
   wire n_19_0_50;
   wire n_19_0_51;
   wire n_19_0_52;
   wire n_19_0_53;
   wire n_19_0_54;
   wire n_19_0_55;
   wire n_19_0_56;
   wire n_19_0_57;
   wire n_19_0_58;
   wire n_19_0_59;
   wire n_19_0_60;
   wire n_19_0_61;
   wire n_19_0_62;
   wire n_19_0_63;
   wire n_19_0_64;
   wire n_19_0_65;
   wire n_19_0_66;
   wire n_19_0_67;
   wire n_19_0_68;
   wire n_19_0_69;
   wire n_19_0_70;
   wire n_19_0_71;
   wire n_19_0_72;
   wire n_19_0_73;
   wire n_19_0_74;
   wire n_19_0_75;
   wire n_19_0_76;
   wire n_19_0_77;
   wire n_19_0_78;
   wire n_19_0_79;
   wire n_19_0_80;
   wire n_19_0_81;
   wire n_19_0_82;
   wire n_19_0_83;
   wire n_19_0_84;
   wire n_19_0_85;
   wire n_19_0_86;
   wire n_19_0_87;
   wire n_19_0_88;
   wire n_19_0_89;
   wire n_19_0_90;
   wire n_19_0_91;
   wire n_19_0_92;
   wire n_19_0_93;
   wire n_19_0_94;
   wire n_19_0_95;
   wire n_19_0_96;
   wire n_19_0_97;
   wire n_19_0_98;
   wire n_19_0_99;
   wire n_19_0_100;
   wire n_19_0_101;
   wire n_19_0_102;
   wire n_19_0_103;
   wire n_19_0_104;
   wire n_19_0_105;
   wire n_19_0_106;
   wire n_19_0_107;
   wire n_19_0_108;
   wire n_19_0_109;
   wire n_19_0_110;
   wire n_19_0_111;
   wire n_19_0_112;
   wire n_19_0_113;
   wire n_19_0_114;
   wire n_19_0_115;
   wire n_19_0_116;
   wire n_19_0_117;
   wire n_19_0_118;
   wire n_19_0_119;
   wire n_19_0_120;
   wire n_19_0_121;
   wire n_19_0_122;
   wire n_19_0_123;
   wire n_19_0_124;
   wire n_19_0_125;
   wire n_19_0_126;
   wire n_19_0_127;
   wire n_19_0_128;
   wire n_19_0_129;
   wire n_19_0_130;
   wire n_19_0_131;
   wire n_19_0_132;
   wire n_19_0_133;
   wire n_19_0_134;
   wire n_19_0_135;
   wire n_19_0_136;
   wire n_19_0_137;
   wire n_19_0_138;
   wire n_19_0_139;
   wire n_19_0_140;
   wire n_19_0_141;
   wire n_19_0_142;
   wire n_19_0_143;
   wire n_19_0_144;
   wire n_19_0_145;
   wire n_19_0_146;
   wire n_19_0_147;
   wire n_19_0_148;
   wire n_19_0_149;
   wire n_19_0_150;
   wire n_19_0_151;
   wire n_19_0_152;
   wire n_19_0_153;
   wire n_19_0_154;
   wire n_19_0_155;
   wire n_19_0_156;
   wire n_19_0_157;
   wire n_19_0_158;
   wire n_19_0_159;
   wire n_19_0_160;
   wire n_19_0_161;
   wire n_19_0_162;
   wire n_19_0_163;
   wire n_19_0_164;
   wire n_19_0_165;
   wire n_19_0_166;
   wire n_19_0_167;

   DFF_X1 \buffer_reg[0][3][3][15]  (.D(\input_filter[3][3] [15]), .CK(n_53_0), 
      .Q(\buffer[0][3][3] [15]), .QN());
   DFF_X1 \buffer_reg[0][3][3][14]  (.D(\input_filter[3][3] [14]), .CK(n_53_0), 
      .Q(\buffer[0][3][3] [14]), .QN());
   DFF_X1 \buffer_reg[0][3][3][13]  (.D(\input_filter[3][3] [13]), .CK(n_53_0), 
      .Q(\buffer[0][3][3] [13]), .QN());
   DFF_X1 \buffer_reg[0][3][3][12]  (.D(\input_filter[3][3] [12]), .CK(n_53_0), 
      .Q(\buffer[0][3][3] [12]), .QN());
   DFF_X1 \buffer_reg[0][3][3][11]  (.D(\input_filter[3][3] [11]), .CK(n_53_0), 
      .Q(\buffer[0][3][3] [11]), .QN());
   DFF_X1 \buffer_reg[0][3][3][10]  (.D(\input_filter[3][3] [10]), .CK(n_53_0), 
      .Q(\buffer[0][3][3] [10]), .QN());
   DFF_X1 \buffer_reg[0][3][3][9]  (.D(\input_filter[3][3] [9]), .CK(n_53_0), 
      .Q(\buffer[0][3][3] [9]), .QN());
   DFF_X1 \buffer_reg[0][3][3][8]  (.D(\input_filter[3][3] [8]), .CK(n_53_0), 
      .Q(\buffer[0][3][3] [8]), .QN());
   DFF_X1 \buffer_reg[0][3][3][7]  (.D(\input_filter[3][3] [7]), .CK(n_53_0), 
      .Q(\buffer[0][3][3] [7]), .QN());
   DFF_X1 \buffer_reg[0][3][3][6]  (.D(\input_filter[3][3] [6]), .CK(n_53_0), 
      .Q(\buffer[0][3][3] [6]), .QN());
   DFF_X1 \buffer_reg[0][3][3][5]  (.D(\input_filter[3][3] [5]), .CK(n_53_0), 
      .Q(\buffer[0][3][3] [5]), .QN());
   DFF_X1 \buffer_reg[0][3][3][4]  (.D(\input_filter[3][3] [4]), .CK(n_53_0), 
      .Q(\buffer[0][3][3] [4]), .QN());
   DFF_X1 \buffer_reg[0][3][3][3]  (.D(\input_filter[3][3] [3]), .CK(n_53_0), 
      .Q(\buffer[0][3][3] [3]), .QN());
   DFF_X1 \buffer_reg[0][3][3][2]  (.D(\input_filter[3][3] [2]), .CK(n_53_0), 
      .Q(\buffer[0][3][3] [2]), .QN());
   DFF_X1 \buffer_reg[0][3][3][1]  (.D(\input_filter[3][3] [1]), .CK(n_53_0), 
      .Q(\buffer[0][3][3] [1]), .QN());
   DFF_X1 \buffer_reg[0][3][3][0]  (.D(\input_filter[3][3] [0]), .CK(n_53_0), 
      .Q(\buffer[0][3][3] [0]), .QN());
   DFF_X1 \buffer_reg[1][3][3][15]  (.D(\input_filter[3][3] [15]), .CK(n_53_1), 
      .Q(\buffer[1][3][3] [15]), .QN());
   DFF_X1 \buffer_reg[1][3][3][14]  (.D(\input_filter[3][3] [14]), .CK(n_53_1), 
      .Q(\buffer[1][3][3] [14]), .QN());
   DFF_X1 \buffer_reg[1][3][3][13]  (.D(\input_filter[3][3] [13]), .CK(n_53_1), 
      .Q(\buffer[1][3][3] [13]), .QN());
   DFF_X1 \buffer_reg[1][3][3][12]  (.D(\input_filter[3][3] [12]), .CK(n_53_1), 
      .Q(\buffer[1][3][3] [12]), .QN());
   DFF_X1 \buffer_reg[1][3][3][11]  (.D(\input_filter[3][3] [11]), .CK(n_53_1), 
      .Q(\buffer[1][3][3] [11]), .QN());
   DFF_X1 \buffer_reg[1][3][3][10]  (.D(\input_filter[3][3] [10]), .CK(n_53_1), 
      .Q(\buffer[1][3][3] [10]), .QN());
   DFF_X1 \buffer_reg[1][3][3][9]  (.D(\input_filter[3][3] [9]), .CK(n_53_1), 
      .Q(\buffer[1][3][3] [9]), .QN());
   DFF_X1 \buffer_reg[1][3][3][8]  (.D(\input_filter[3][3] [8]), .CK(n_53_1), 
      .Q(\buffer[1][3][3] [8]), .QN());
   DFF_X1 \buffer_reg[1][3][3][7]  (.D(\input_filter[3][3] [7]), .CK(n_53_1), 
      .Q(\buffer[1][3][3] [7]), .QN());
   DFF_X1 \buffer_reg[1][3][3][6]  (.D(\input_filter[3][3] [6]), .CK(n_53_1), 
      .Q(\buffer[1][3][3] [6]), .QN());
   DFF_X1 \buffer_reg[1][3][3][5]  (.D(\input_filter[3][3] [5]), .CK(n_53_1), 
      .Q(\buffer[1][3][3] [5]), .QN());
   DFF_X1 \buffer_reg[1][3][3][4]  (.D(\input_filter[3][3] [4]), .CK(n_53_1), 
      .Q(\buffer[1][3][3] [4]), .QN());
   DFF_X1 \buffer_reg[1][3][3][3]  (.D(\input_filter[3][3] [3]), .CK(n_53_1), 
      .Q(\buffer[1][3][3] [3]), .QN());
   DFF_X1 \buffer_reg[1][3][3][2]  (.D(\input_filter[3][3] [2]), .CK(n_53_1), 
      .Q(\buffer[1][3][3] [2]), .QN());
   DFF_X1 \buffer_reg[1][3][3][1]  (.D(\input_filter[3][3] [1]), .CK(n_53_1), 
      .Q(\buffer[1][3][3] [1]), .QN());
   DFF_X1 \buffer_reg[1][3][3][0]  (.D(\input_filter[3][3] [0]), .CK(n_53_1), 
      .Q(\buffer[1][3][3] [0]), .QN());
   DFF_X1 \buffer_reg[2][3][3][15]  (.D(\input_filter[3][3] [15]), .CK(n_53_2), 
      .Q(\buffer[2][3][3] [15]), .QN());
   DFF_X1 \buffer_reg[2][3][3][14]  (.D(\input_filter[3][3] [14]), .CK(n_53_2), 
      .Q(\buffer[2][3][3] [14]), .QN());
   DFF_X1 \buffer_reg[2][3][3][13]  (.D(\input_filter[3][3] [13]), .CK(n_53_2), 
      .Q(\buffer[2][3][3] [13]), .QN());
   DFF_X1 \buffer_reg[2][3][3][12]  (.D(\input_filter[3][3] [12]), .CK(n_53_2), 
      .Q(\buffer[2][3][3] [12]), .QN());
   DFF_X1 \buffer_reg[2][3][3][11]  (.D(\input_filter[3][3] [11]), .CK(n_53_2), 
      .Q(\buffer[2][3][3] [11]), .QN());
   DFF_X1 \buffer_reg[2][3][3][10]  (.D(\input_filter[3][3] [10]), .CK(n_53_2), 
      .Q(\buffer[2][3][3] [10]), .QN());
   DFF_X1 \buffer_reg[2][3][3][9]  (.D(\input_filter[3][3] [9]), .CK(n_53_2), 
      .Q(\buffer[2][3][3] [9]), .QN());
   DFF_X1 \buffer_reg[2][3][3][8]  (.D(\input_filter[3][3] [8]), .CK(n_53_2), 
      .Q(\buffer[2][3][3] [8]), .QN());
   DFF_X1 \buffer_reg[2][3][3][7]  (.D(\input_filter[3][3] [7]), .CK(n_53_2), 
      .Q(\buffer[2][3][3] [7]), .QN());
   DFF_X1 \buffer_reg[2][3][3][6]  (.D(\input_filter[3][3] [6]), .CK(n_53_2), 
      .Q(\buffer[2][3][3] [6]), .QN());
   DFF_X1 \buffer_reg[2][3][3][5]  (.D(\input_filter[3][3] [5]), .CK(n_53_2), 
      .Q(\buffer[2][3][3] [5]), .QN());
   DFF_X1 \buffer_reg[2][3][3][4]  (.D(\input_filter[3][3] [4]), .CK(n_53_2), 
      .Q(\buffer[2][3][3] [4]), .QN());
   DFF_X1 \buffer_reg[2][3][3][3]  (.D(\input_filter[3][3] [3]), .CK(n_53_2), 
      .Q(\buffer[2][3][3] [3]), .QN());
   DFF_X1 \buffer_reg[2][3][3][2]  (.D(\input_filter[3][3] [2]), .CK(n_53_2), 
      .Q(\buffer[2][3][3] [2]), .QN());
   DFF_X1 \buffer_reg[2][3][3][1]  (.D(\input_filter[3][3] [1]), .CK(n_53_2), 
      .Q(\buffer[2][3][3] [1]), .QN());
   DFF_X1 \buffer_reg[2][3][3][0]  (.D(\input_filter[3][3] [0]), .CK(n_53_2), 
      .Q(\buffer[2][3][3] [0]), .QN());
   DFF_X1 \buffer_reg[3][3][3][15]  (.D(\input_filter[3][3] [15]), .CK(n_53_3), 
      .Q(\buffer[3][3][3] [15]), .QN());
   DFF_X1 \buffer_reg[3][3][3][14]  (.D(\input_filter[3][3] [14]), .CK(n_53_3), 
      .Q(\buffer[3][3][3] [14]), .QN());
   DFF_X1 \buffer_reg[3][3][3][13]  (.D(\input_filter[3][3] [13]), .CK(n_53_3), 
      .Q(\buffer[3][3][3] [13]), .QN());
   DFF_X1 \buffer_reg[3][3][3][12]  (.D(\input_filter[3][3] [12]), .CK(n_53_3), 
      .Q(\buffer[3][3][3] [12]), .QN());
   DFF_X1 \buffer_reg[3][3][3][11]  (.D(\input_filter[3][3] [11]), .CK(n_53_3), 
      .Q(\buffer[3][3][3] [11]), .QN());
   DFF_X1 \buffer_reg[3][3][3][10]  (.D(\input_filter[3][3] [10]), .CK(n_53_3), 
      .Q(\buffer[3][3][3] [10]), .QN());
   DFF_X1 \buffer_reg[3][3][3][9]  (.D(\input_filter[3][3] [9]), .CK(n_53_3), 
      .Q(\buffer[3][3][3] [9]), .QN());
   DFF_X1 \buffer_reg[3][3][3][8]  (.D(\input_filter[3][3] [8]), .CK(n_53_3), 
      .Q(\buffer[3][3][3] [8]), .QN());
   DFF_X1 \buffer_reg[3][3][3][7]  (.D(\input_filter[3][3] [7]), .CK(n_53_3), 
      .Q(\buffer[3][3][3] [7]), .QN());
   DFF_X1 \buffer_reg[3][3][3][6]  (.D(\input_filter[3][3] [6]), .CK(n_53_3), 
      .Q(\buffer[3][3][3] [6]), .QN());
   DFF_X1 \buffer_reg[3][3][3][5]  (.D(\input_filter[3][3] [5]), .CK(n_53_3), 
      .Q(\buffer[3][3][3] [5]), .QN());
   DFF_X1 \buffer_reg[3][3][3][4]  (.D(\input_filter[3][3] [4]), .CK(n_53_3), 
      .Q(\buffer[3][3][3] [4]), .QN());
   DFF_X1 \buffer_reg[3][3][3][3]  (.D(\input_filter[3][3] [3]), .CK(n_53_3), 
      .Q(\buffer[3][3][3] [3]), .QN());
   DFF_X1 \buffer_reg[3][3][3][2]  (.D(\input_filter[3][3] [2]), .CK(n_53_3), 
      .Q(\buffer[3][3][3] [2]), .QN());
   DFF_X1 \buffer_reg[3][3][3][1]  (.D(\input_filter[3][3] [1]), .CK(n_53_3), 
      .Q(\buffer[3][3][3] [1]), .QN());
   DFF_X1 \buffer_reg[3][3][3][0]  (.D(\input_filter[3][3] [0]), .CK(n_53_3), 
      .Q(\buffer[3][3][3] [0]), .QN());
   DFF_X1 \buffer_reg[4][3][3][15]  (.D(\input_filter[3][3] [15]), .CK(n_53_4), 
      .Q(\buffer[4][3][3] [15]), .QN());
   DFF_X1 \buffer_reg[4][3][3][14]  (.D(\input_filter[3][3] [14]), .CK(n_53_4), 
      .Q(\buffer[4][3][3] [14]), .QN());
   DFF_X1 \buffer_reg[4][3][3][13]  (.D(\input_filter[3][3] [13]), .CK(n_53_4), 
      .Q(\buffer[4][3][3] [13]), .QN());
   DFF_X1 \buffer_reg[4][3][3][12]  (.D(\input_filter[3][3] [12]), .CK(n_53_4), 
      .Q(\buffer[4][3][3] [12]), .QN());
   DFF_X1 \buffer_reg[4][3][3][11]  (.D(\input_filter[3][3] [11]), .CK(n_53_4), 
      .Q(\buffer[4][3][3] [11]), .QN());
   DFF_X1 \buffer_reg[4][3][3][10]  (.D(\input_filter[3][3] [10]), .CK(n_53_4), 
      .Q(\buffer[4][3][3] [10]), .QN());
   DFF_X1 \buffer_reg[4][3][3][9]  (.D(\input_filter[3][3] [9]), .CK(n_53_4), 
      .Q(\buffer[4][3][3] [9]), .QN());
   DFF_X1 \buffer_reg[4][3][3][8]  (.D(\input_filter[3][3] [8]), .CK(n_53_4), 
      .Q(\buffer[4][3][3] [8]), .QN());
   DFF_X1 \buffer_reg[4][3][3][7]  (.D(\input_filter[3][3] [7]), .CK(n_53_4), 
      .Q(\buffer[4][3][3] [7]), .QN());
   DFF_X1 \buffer_reg[4][3][3][6]  (.D(\input_filter[3][3] [6]), .CK(n_53_4), 
      .Q(\buffer[4][3][3] [6]), .QN());
   DFF_X1 \buffer_reg[4][3][3][5]  (.D(\input_filter[3][3] [5]), .CK(n_53_4), 
      .Q(\buffer[4][3][3] [5]), .QN());
   DFF_X1 \buffer_reg[4][3][3][4]  (.D(\input_filter[3][3] [4]), .CK(n_53_4), 
      .Q(\buffer[4][3][3] [4]), .QN());
   DFF_X1 \buffer_reg[4][3][3][3]  (.D(\input_filter[3][3] [3]), .CK(n_53_4), 
      .Q(\buffer[4][3][3] [3]), .QN());
   DFF_X1 \buffer_reg[4][3][3][2]  (.D(\input_filter[3][3] [2]), .CK(n_53_4), 
      .Q(\buffer[4][3][3] [2]), .QN());
   DFF_X1 \buffer_reg[4][3][3][1]  (.D(\input_filter[3][3] [1]), .CK(n_53_4), 
      .Q(\buffer[4][3][3] [1]), .QN());
   DFF_X1 \buffer_reg[4][3][3][0]  (.D(\input_filter[3][3] [0]), .CK(n_53_4), 
      .Q(\buffer[4][3][3] [0]), .QN());
   DFF_X1 \buffer_reg[5][3][3][15]  (.D(\input_filter[3][3] [15]), .CK(n_53_5), 
      .Q(\buffer[5][3][3] [15]), .QN());
   DFF_X1 \buffer_reg[5][3][3][14]  (.D(\input_filter[3][3] [14]), .CK(n_53_5), 
      .Q(\buffer[5][3][3] [14]), .QN());
   DFF_X1 \buffer_reg[5][3][3][13]  (.D(\input_filter[3][3] [13]), .CK(n_53_5), 
      .Q(\buffer[5][3][3] [13]), .QN());
   DFF_X1 \buffer_reg[5][3][3][12]  (.D(\input_filter[3][3] [12]), .CK(n_53_5), 
      .Q(\buffer[5][3][3] [12]), .QN());
   DFF_X1 \buffer_reg[5][3][3][11]  (.D(\input_filter[3][3] [11]), .CK(n_53_5), 
      .Q(\buffer[5][3][3] [11]), .QN());
   DFF_X1 \buffer_reg[5][3][3][10]  (.D(\input_filter[3][3] [10]), .CK(n_53_5), 
      .Q(\buffer[5][3][3] [10]), .QN());
   DFF_X1 \buffer_reg[5][3][3][9]  (.D(\input_filter[3][3] [9]), .CK(n_53_5), 
      .Q(\buffer[5][3][3] [9]), .QN());
   DFF_X1 \buffer_reg[5][3][3][8]  (.D(\input_filter[3][3] [8]), .CK(n_53_5), 
      .Q(\buffer[5][3][3] [8]), .QN());
   DFF_X1 \buffer_reg[5][3][3][7]  (.D(\input_filter[3][3] [7]), .CK(n_53_5), 
      .Q(\buffer[5][3][3] [7]), .QN());
   DFF_X1 \buffer_reg[5][3][3][6]  (.D(\input_filter[3][3] [6]), .CK(n_53_5), 
      .Q(\buffer[5][3][3] [6]), .QN());
   DFF_X1 \buffer_reg[5][3][3][5]  (.D(\input_filter[3][3] [5]), .CK(n_53_5), 
      .Q(\buffer[5][3][3] [5]), .QN());
   DFF_X1 \buffer_reg[5][3][3][4]  (.D(\input_filter[3][3] [4]), .CK(n_53_5), 
      .Q(\buffer[5][3][3] [4]), .QN());
   DFF_X1 \buffer_reg[5][3][3][3]  (.D(\input_filter[3][3] [3]), .CK(n_53_5), 
      .Q(\buffer[5][3][3] [3]), .QN());
   DFF_X1 \buffer_reg[5][3][3][2]  (.D(\input_filter[3][3] [2]), .CK(n_53_5), 
      .Q(\buffer[5][3][3] [2]), .QN());
   DFF_X1 \buffer_reg[5][3][3][1]  (.D(\input_filter[3][3] [1]), .CK(n_53_5), 
      .Q(\buffer[5][3][3] [1]), .QN());
   DFF_X1 \buffer_reg[5][3][3][0]  (.D(\input_filter[3][3] [0]), .CK(n_53_5), 
      .Q(\buffer[5][3][3] [0]), .QN());
   DFF_X1 \buffer_reg[6][3][3][15]  (.D(\input_filter[3][3] [15]), .CK(n_53_6), 
      .Q(\buffer[6][3][3] [15]), .QN());
   DFF_X1 \buffer_reg[6][3][3][14]  (.D(\input_filter[3][3] [14]), .CK(n_53_6), 
      .Q(\buffer[6][3][3] [14]), .QN());
   DFF_X1 \buffer_reg[6][3][3][13]  (.D(\input_filter[3][3] [13]), .CK(n_53_6), 
      .Q(\buffer[6][3][3] [13]), .QN());
   DFF_X1 \buffer_reg[6][3][3][12]  (.D(\input_filter[3][3] [12]), .CK(n_53_6), 
      .Q(\buffer[6][3][3] [12]), .QN());
   DFF_X1 \buffer_reg[6][3][3][11]  (.D(\input_filter[3][3] [11]), .CK(n_53_6), 
      .Q(\buffer[6][3][3] [11]), .QN());
   DFF_X1 \buffer_reg[6][3][3][10]  (.D(\input_filter[3][3] [10]), .CK(n_53_6), 
      .Q(\buffer[6][3][3] [10]), .QN());
   DFF_X1 \buffer_reg[6][3][3][9]  (.D(\input_filter[3][3] [9]), .CK(n_53_6), 
      .Q(\buffer[6][3][3] [9]), .QN());
   DFF_X1 \buffer_reg[6][3][3][8]  (.D(\input_filter[3][3] [8]), .CK(n_53_6), 
      .Q(\buffer[6][3][3] [8]), .QN());
   DFF_X1 \buffer_reg[6][3][3][7]  (.D(\input_filter[3][3] [7]), .CK(n_53_6), 
      .Q(\buffer[6][3][3] [7]), .QN());
   DFF_X1 \buffer_reg[6][3][3][6]  (.D(\input_filter[3][3] [6]), .CK(n_53_6), 
      .Q(\buffer[6][3][3] [6]), .QN());
   DFF_X1 \buffer_reg[6][3][3][5]  (.D(\input_filter[3][3] [5]), .CK(n_53_6), 
      .Q(\buffer[6][3][3] [5]), .QN());
   DFF_X1 \buffer_reg[6][3][3][4]  (.D(\input_filter[3][3] [4]), .CK(n_53_6), 
      .Q(\buffer[6][3][3] [4]), .QN());
   DFF_X1 \buffer_reg[6][3][3][3]  (.D(\input_filter[3][3] [3]), .CK(n_53_6), 
      .Q(\buffer[6][3][3] [3]), .QN());
   DFF_X1 \buffer_reg[6][3][3][2]  (.D(\input_filter[3][3] [2]), .CK(n_53_6), 
      .Q(\buffer[6][3][3] [2]), .QN());
   DFF_X1 \buffer_reg[6][3][3][1]  (.D(\input_filter[3][3] [1]), .CK(n_53_6), 
      .Q(\buffer[6][3][3] [1]), .QN());
   DFF_X1 \buffer_reg[6][3][3][0]  (.D(\input_filter[3][3] [0]), .CK(n_53_6), 
      .Q(\buffer[6][3][3] [0]), .QN());
   DFF_X1 \buffer_reg[7][3][3][15]  (.D(\input_filter[3][3] [15]), .CK(n_53_7), 
      .Q(\buffer[7][3][3] [15]), .QN());
   DFF_X1 \buffer_reg[7][3][3][14]  (.D(\input_filter[3][3] [14]), .CK(n_53_7), 
      .Q(\buffer[7][3][3] [14]), .QN());
   DFF_X1 \buffer_reg[7][3][3][13]  (.D(\input_filter[3][3] [13]), .CK(n_53_7), 
      .Q(\buffer[7][3][3] [13]), .QN());
   DFF_X1 \buffer_reg[7][3][3][12]  (.D(\input_filter[3][3] [12]), .CK(n_53_7), 
      .Q(\buffer[7][3][3] [12]), .QN());
   DFF_X1 \buffer_reg[7][3][3][11]  (.D(\input_filter[3][3] [11]), .CK(n_53_7), 
      .Q(\buffer[7][3][3] [11]), .QN());
   DFF_X1 \buffer_reg[7][3][3][10]  (.D(\input_filter[3][3] [10]), .CK(n_53_7), 
      .Q(\buffer[7][3][3] [10]), .QN());
   DFF_X1 \buffer_reg[7][3][3][9]  (.D(\input_filter[3][3] [9]), .CK(n_53_7), 
      .Q(\buffer[7][3][3] [9]), .QN());
   DFF_X1 \buffer_reg[7][3][3][8]  (.D(\input_filter[3][3] [8]), .CK(n_53_7), 
      .Q(\buffer[7][3][3] [8]), .QN());
   DFF_X1 \buffer_reg[7][3][3][7]  (.D(\input_filter[3][3] [7]), .CK(n_53_7), 
      .Q(\buffer[7][3][3] [7]), .QN());
   DFF_X1 \buffer_reg[7][3][3][6]  (.D(\input_filter[3][3] [6]), .CK(n_53_7), 
      .Q(\buffer[7][3][3] [6]), .QN());
   DFF_X1 \buffer_reg[7][3][3][5]  (.D(\input_filter[3][3] [5]), .CK(n_53_7), 
      .Q(\buffer[7][3][3] [5]), .QN());
   DFF_X1 \buffer_reg[7][3][3][4]  (.D(\input_filter[3][3] [4]), .CK(n_53_7), 
      .Q(\buffer[7][3][3] [4]), .QN());
   DFF_X1 \buffer_reg[7][3][3][3]  (.D(\input_filter[3][3] [3]), .CK(n_53_7), 
      .Q(\buffer[7][3][3] [3]), .QN());
   DFF_X1 \buffer_reg[7][3][3][2]  (.D(\input_filter[3][3] [2]), .CK(n_53_7), 
      .Q(\buffer[7][3][3] [2]), .QN());
   DFF_X1 \buffer_reg[7][3][3][1]  (.D(\input_filter[3][3] [1]), .CK(n_53_7), 
      .Q(\buffer[7][3][3] [1]), .QN());
   DFF_X1 \buffer_reg[7][3][3][0]  (.D(\input_filter[3][3] [0]), .CK(n_53_7), 
      .Q(\buffer[7][3][3] [0]), .QN());
   DFF_X1 \buffer_reg[8][3][3][15]  (.D(\input_filter[3][3] [15]), .CK(n_53_8), 
      .Q(\buffer[8][3][3] [15]), .QN());
   DFF_X1 \buffer_reg[8][3][3][14]  (.D(\input_filter[3][3] [14]), .CK(n_53_8), 
      .Q(\buffer[8][3][3] [14]), .QN());
   DFF_X1 \buffer_reg[8][3][3][13]  (.D(\input_filter[3][3] [13]), .CK(n_53_8), 
      .Q(\buffer[8][3][3] [13]), .QN());
   DFF_X1 \buffer_reg[8][3][3][12]  (.D(\input_filter[3][3] [12]), .CK(n_53_8), 
      .Q(\buffer[8][3][3] [12]), .QN());
   DFF_X1 \buffer_reg[8][3][3][11]  (.D(\input_filter[3][3] [11]), .CK(n_53_8), 
      .Q(\buffer[8][3][3] [11]), .QN());
   DFF_X1 \buffer_reg[8][3][3][10]  (.D(\input_filter[3][3] [10]), .CK(n_53_8), 
      .Q(\buffer[8][3][3] [10]), .QN());
   DFF_X1 \buffer_reg[8][3][3][9]  (.D(\input_filter[3][3] [9]), .CK(n_53_8), 
      .Q(\buffer[8][3][3] [9]), .QN());
   DFF_X1 \buffer_reg[8][3][3][8]  (.D(\input_filter[3][3] [8]), .CK(n_53_8), 
      .Q(\buffer[8][3][3] [8]), .QN());
   DFF_X1 \buffer_reg[8][3][3][7]  (.D(\input_filter[3][3] [7]), .CK(n_53_8), 
      .Q(\buffer[8][3][3] [7]), .QN());
   DFF_X1 \buffer_reg[8][3][3][6]  (.D(\input_filter[3][3] [6]), .CK(n_53_8), 
      .Q(\buffer[8][3][3] [6]), .QN());
   DFF_X1 \buffer_reg[8][3][3][5]  (.D(\input_filter[3][3] [5]), .CK(n_53_8), 
      .Q(\buffer[8][3][3] [5]), .QN());
   DFF_X1 \buffer_reg[8][3][3][4]  (.D(\input_filter[3][3] [4]), .CK(n_53_8), 
      .Q(\buffer[8][3][3] [4]), .QN());
   DFF_X1 \buffer_reg[8][3][3][3]  (.D(\input_filter[3][3] [3]), .CK(n_53_8), 
      .Q(\buffer[8][3][3] [3]), .QN());
   DFF_X1 \buffer_reg[8][3][3][2]  (.D(\input_filter[3][3] [2]), .CK(n_53_8), 
      .Q(\buffer[8][3][3] [2]), .QN());
   DFF_X1 \buffer_reg[8][3][3][1]  (.D(\input_filter[3][3] [1]), .CK(n_53_8), 
      .Q(\buffer[8][3][3] [1]), .QN());
   DFF_X1 \buffer_reg[8][3][3][0]  (.D(\input_filter[3][3] [0]), .CK(n_53_8), 
      .Q(\buffer[8][3][3] [0]), .QN());
   DFF_X1 \buffer_reg[9][3][3][15]  (.D(\input_filter[3][3] [15]), .CK(n_53_9), 
      .Q(\buffer[9][3][3] [15]), .QN());
   DFF_X1 \buffer_reg[9][3][3][14]  (.D(\input_filter[3][3] [14]), .CK(n_53_9), 
      .Q(\buffer[9][3][3] [14]), .QN());
   DFF_X1 \buffer_reg[9][3][3][13]  (.D(\input_filter[3][3] [13]), .CK(n_53_9), 
      .Q(\buffer[9][3][3] [13]), .QN());
   DFF_X1 \buffer_reg[9][3][3][12]  (.D(\input_filter[3][3] [12]), .CK(n_53_9), 
      .Q(\buffer[9][3][3] [12]), .QN());
   DFF_X1 \buffer_reg[9][3][3][11]  (.D(\input_filter[3][3] [11]), .CK(n_53_9), 
      .Q(\buffer[9][3][3] [11]), .QN());
   DFF_X1 \buffer_reg[9][3][3][10]  (.D(\input_filter[3][3] [10]), .CK(n_53_9), 
      .Q(\buffer[9][3][3] [10]), .QN());
   DFF_X1 \buffer_reg[9][3][3][9]  (.D(\input_filter[3][3] [9]), .CK(n_53_9), 
      .Q(\buffer[9][3][3] [9]), .QN());
   DFF_X1 \buffer_reg[9][3][3][8]  (.D(\input_filter[3][3] [8]), .CK(n_53_9), 
      .Q(\buffer[9][3][3] [8]), .QN());
   DFF_X1 \buffer_reg[9][3][3][7]  (.D(\input_filter[3][3] [7]), .CK(n_53_9), 
      .Q(\buffer[9][3][3] [7]), .QN());
   DFF_X1 \buffer_reg[9][3][3][6]  (.D(\input_filter[3][3] [6]), .CK(n_53_9), 
      .Q(\buffer[9][3][3] [6]), .QN());
   DFF_X1 \buffer_reg[9][3][3][5]  (.D(\input_filter[3][3] [5]), .CK(n_53_9), 
      .Q(\buffer[9][3][3] [5]), .QN());
   DFF_X1 \buffer_reg[9][3][3][4]  (.D(\input_filter[3][3] [4]), .CK(n_53_9), 
      .Q(\buffer[9][3][3] [4]), .QN());
   DFF_X1 \buffer_reg[9][3][3][3]  (.D(\input_filter[3][3] [3]), .CK(n_53_9), 
      .Q(\buffer[9][3][3] [3]), .QN());
   DFF_X1 \buffer_reg[9][3][3][2]  (.D(\input_filter[3][3] [2]), .CK(n_53_9), 
      .Q(\buffer[9][3][3] [2]), .QN());
   DFF_X1 \buffer_reg[9][3][3][1]  (.D(\input_filter[3][3] [1]), .CK(n_53_9), 
      .Q(\buffer[9][3][3] [1]), .QN());
   DFF_X1 \buffer_reg[9][3][3][0]  (.D(\input_filter[3][3] [0]), .CK(n_53_9), 
      .Q(\buffer[9][3][3] [0]), .QN());
   DFF_X1 \buffer_reg[10][3][3][15]  (.D(\input_filter[3][3] [15]), .CK(n_53_10), 
      .Q(\buffer[10][3][3] [15]), .QN());
   DFF_X1 \buffer_reg[10][3][3][14]  (.D(\input_filter[3][3] [14]), .CK(n_53_10), 
      .Q(\buffer[10][3][3] [14]), .QN());
   DFF_X1 \buffer_reg[10][3][3][13]  (.D(\input_filter[3][3] [13]), .CK(n_53_10), 
      .Q(\buffer[10][3][3] [13]), .QN());
   DFF_X1 \buffer_reg[10][3][3][12]  (.D(\input_filter[3][3] [12]), .CK(n_53_10), 
      .Q(\buffer[10][3][3] [12]), .QN());
   DFF_X1 \buffer_reg[10][3][3][11]  (.D(\input_filter[3][3] [11]), .CK(n_53_10), 
      .Q(\buffer[10][3][3] [11]), .QN());
   DFF_X1 \buffer_reg[10][3][3][10]  (.D(\input_filter[3][3] [10]), .CK(n_53_10), 
      .Q(\buffer[10][3][3] [10]), .QN());
   DFF_X1 \buffer_reg[10][3][3][9]  (.D(\input_filter[3][3] [9]), .CK(n_53_10), 
      .Q(\buffer[10][3][3] [9]), .QN());
   DFF_X1 \buffer_reg[10][3][3][8]  (.D(\input_filter[3][3] [8]), .CK(n_53_10), 
      .Q(\buffer[10][3][3] [8]), .QN());
   DFF_X1 \buffer_reg[10][3][3][7]  (.D(\input_filter[3][3] [7]), .CK(n_53_10), 
      .Q(\buffer[10][3][3] [7]), .QN());
   DFF_X1 \buffer_reg[10][3][3][6]  (.D(\input_filter[3][3] [6]), .CK(n_53_10), 
      .Q(\buffer[10][3][3] [6]), .QN());
   DFF_X1 \buffer_reg[10][3][3][5]  (.D(\input_filter[3][3] [5]), .CK(n_53_10), 
      .Q(\buffer[10][3][3] [5]), .QN());
   DFF_X1 \buffer_reg[10][3][3][4]  (.D(\input_filter[3][3] [4]), .CK(n_53_10), 
      .Q(\buffer[10][3][3] [4]), .QN());
   DFF_X1 \buffer_reg[10][3][3][3]  (.D(\input_filter[3][3] [3]), .CK(n_53_10), 
      .Q(\buffer[10][3][3] [3]), .QN());
   DFF_X1 \buffer_reg[10][3][3][2]  (.D(\input_filter[3][3] [2]), .CK(n_53_10), 
      .Q(\buffer[10][3][3] [2]), .QN());
   DFF_X1 \buffer_reg[10][3][3][1]  (.D(\input_filter[3][3] [1]), .CK(n_53_10), 
      .Q(\buffer[10][3][3] [1]), .QN());
   DFF_X1 \buffer_reg[10][3][3][0]  (.D(\input_filter[3][3] [0]), .CK(n_53_10), 
      .Q(\buffer[10][3][3] [0]), .QN());
   DFF_X1 \buffer_reg[11][3][3][15]  (.D(\input_filter[3][3] [15]), .CK(n_53_11), 
      .Q(\buffer[11][3][3] [15]), .QN());
   DFF_X1 \buffer_reg[11][3][3][14]  (.D(\input_filter[3][3] [14]), .CK(n_53_11), 
      .Q(\buffer[11][3][3] [14]), .QN());
   DFF_X1 \buffer_reg[11][3][3][13]  (.D(\input_filter[3][3] [13]), .CK(n_53_11), 
      .Q(\buffer[11][3][3] [13]), .QN());
   DFF_X1 \buffer_reg[11][3][3][12]  (.D(\input_filter[3][3] [12]), .CK(n_53_11), 
      .Q(\buffer[11][3][3] [12]), .QN());
   DFF_X1 \buffer_reg[11][3][3][11]  (.D(\input_filter[3][3] [11]), .CK(n_53_11), 
      .Q(\buffer[11][3][3] [11]), .QN());
   DFF_X1 \buffer_reg[11][3][3][10]  (.D(\input_filter[3][3] [10]), .CK(n_53_11), 
      .Q(\buffer[11][3][3] [10]), .QN());
   DFF_X1 \buffer_reg[11][3][3][9]  (.D(\input_filter[3][3] [9]), .CK(n_53_11), 
      .Q(\buffer[11][3][3] [9]), .QN());
   DFF_X1 \buffer_reg[11][3][3][8]  (.D(\input_filter[3][3] [8]), .CK(n_53_11), 
      .Q(\buffer[11][3][3] [8]), .QN());
   DFF_X1 \buffer_reg[11][3][3][7]  (.D(\input_filter[3][3] [7]), .CK(n_53_11), 
      .Q(\buffer[11][3][3] [7]), .QN());
   DFF_X1 \buffer_reg[11][3][3][6]  (.D(\input_filter[3][3] [6]), .CK(n_53_11), 
      .Q(\buffer[11][3][3] [6]), .QN());
   DFF_X1 \buffer_reg[11][3][3][5]  (.D(\input_filter[3][3] [5]), .CK(n_53_11), 
      .Q(\buffer[11][3][3] [5]), .QN());
   DFF_X1 \buffer_reg[11][3][3][4]  (.D(\input_filter[3][3] [4]), .CK(n_53_11), 
      .Q(\buffer[11][3][3] [4]), .QN());
   DFF_X1 \buffer_reg[11][3][3][3]  (.D(\input_filter[3][3] [3]), .CK(n_53_11), 
      .Q(\buffer[11][3][3] [3]), .QN());
   DFF_X1 \buffer_reg[11][3][3][2]  (.D(\input_filter[3][3] [2]), .CK(n_53_11), 
      .Q(\buffer[11][3][3] [2]), .QN());
   DFF_X1 \buffer_reg[11][3][3][1]  (.D(\input_filter[3][3] [1]), .CK(n_53_11), 
      .Q(\buffer[11][3][3] [1]), .QN());
   DFF_X1 \buffer_reg[11][3][3][0]  (.D(\input_filter[3][3] [0]), .CK(n_53_11), 
      .Q(\buffer[11][3][3] [0]), .QN());
   DFF_X1 \buffer_reg[12][3][3][15]  (.D(\input_filter[3][3] [15]), .CK(n_53_12), 
      .Q(\buffer[12][3][3] [15]), .QN());
   DFF_X1 \buffer_reg[12][3][3][14]  (.D(\input_filter[3][3] [14]), .CK(n_53_12), 
      .Q(\buffer[12][3][3] [14]), .QN());
   DFF_X1 \buffer_reg[12][3][3][13]  (.D(\input_filter[3][3] [13]), .CK(n_53_12), 
      .Q(\buffer[12][3][3] [13]), .QN());
   DFF_X1 \buffer_reg[12][3][3][12]  (.D(\input_filter[3][3] [12]), .CK(n_53_12), 
      .Q(\buffer[12][3][3] [12]), .QN());
   DFF_X1 \buffer_reg[12][3][3][11]  (.D(\input_filter[3][3] [11]), .CK(n_53_12), 
      .Q(\buffer[12][3][3] [11]), .QN());
   DFF_X1 \buffer_reg[12][3][3][10]  (.D(\input_filter[3][3] [10]), .CK(n_53_12), 
      .Q(\buffer[12][3][3] [10]), .QN());
   DFF_X1 \buffer_reg[12][3][3][9]  (.D(\input_filter[3][3] [9]), .CK(n_53_12), 
      .Q(\buffer[12][3][3] [9]), .QN());
   DFF_X1 \buffer_reg[12][3][3][8]  (.D(\input_filter[3][3] [8]), .CK(n_53_12), 
      .Q(\buffer[12][3][3] [8]), .QN());
   DFF_X1 \buffer_reg[12][3][3][7]  (.D(\input_filter[3][3] [7]), .CK(n_53_12), 
      .Q(\buffer[12][3][3] [7]), .QN());
   DFF_X1 \buffer_reg[12][3][3][6]  (.D(\input_filter[3][3] [6]), .CK(n_53_12), 
      .Q(\buffer[12][3][3] [6]), .QN());
   DFF_X1 \buffer_reg[12][3][3][5]  (.D(\input_filter[3][3] [5]), .CK(n_53_12), 
      .Q(\buffer[12][3][3] [5]), .QN());
   DFF_X1 \buffer_reg[12][3][3][4]  (.D(\input_filter[3][3] [4]), .CK(n_53_12), 
      .Q(\buffer[12][3][3] [4]), .QN());
   DFF_X1 \buffer_reg[12][3][3][3]  (.D(\input_filter[3][3] [3]), .CK(n_53_12), 
      .Q(\buffer[12][3][3] [3]), .QN());
   DFF_X1 \buffer_reg[12][3][3][2]  (.D(\input_filter[3][3] [2]), .CK(n_53_12), 
      .Q(\buffer[12][3][3] [2]), .QN());
   DFF_X1 \buffer_reg[12][3][3][1]  (.D(\input_filter[3][3] [1]), .CK(n_53_12), 
      .Q(\buffer[12][3][3] [1]), .QN());
   DFF_X1 \buffer_reg[12][3][3][0]  (.D(\input_filter[3][3] [0]), .CK(n_53_12), 
      .Q(\buffer[12][3][3] [0]), .QN());
   DFF_X1 \buffer_reg[13][3][3][15]  (.D(\input_filter[3][3] [15]), .CK(n_53_13), 
      .Q(\buffer[13][3][3] [15]), .QN());
   DFF_X1 \buffer_reg[13][3][3][14]  (.D(\input_filter[3][3] [14]), .CK(n_53_13), 
      .Q(\buffer[13][3][3] [14]), .QN());
   DFF_X1 \buffer_reg[13][3][3][13]  (.D(\input_filter[3][3] [13]), .CK(n_53_13), 
      .Q(\buffer[13][3][3] [13]), .QN());
   DFF_X1 \buffer_reg[13][3][3][12]  (.D(\input_filter[3][3] [12]), .CK(n_53_13), 
      .Q(\buffer[13][3][3] [12]), .QN());
   DFF_X1 \buffer_reg[13][3][3][11]  (.D(\input_filter[3][3] [11]), .CK(n_53_13), 
      .Q(\buffer[13][3][3] [11]), .QN());
   DFF_X1 \buffer_reg[13][3][3][10]  (.D(\input_filter[3][3] [10]), .CK(n_53_13), 
      .Q(\buffer[13][3][3] [10]), .QN());
   DFF_X1 \buffer_reg[13][3][3][9]  (.D(\input_filter[3][3] [9]), .CK(n_53_13), 
      .Q(\buffer[13][3][3] [9]), .QN());
   DFF_X1 \buffer_reg[13][3][3][8]  (.D(\input_filter[3][3] [8]), .CK(n_53_13), 
      .Q(\buffer[13][3][3] [8]), .QN());
   DFF_X1 \buffer_reg[13][3][3][7]  (.D(\input_filter[3][3] [7]), .CK(n_53_13), 
      .Q(\buffer[13][3][3] [7]), .QN());
   DFF_X1 \buffer_reg[13][3][3][6]  (.D(\input_filter[3][3] [6]), .CK(n_53_13), 
      .Q(\buffer[13][3][3] [6]), .QN());
   DFF_X1 \buffer_reg[13][3][3][5]  (.D(\input_filter[3][3] [5]), .CK(n_53_13), 
      .Q(\buffer[13][3][3] [5]), .QN());
   DFF_X1 \buffer_reg[13][3][3][4]  (.D(\input_filter[3][3] [4]), .CK(n_53_13), 
      .Q(\buffer[13][3][3] [4]), .QN());
   DFF_X1 \buffer_reg[13][3][3][3]  (.D(\input_filter[3][3] [3]), .CK(n_53_13), 
      .Q(\buffer[13][3][3] [3]), .QN());
   DFF_X1 \buffer_reg[13][3][3][2]  (.D(\input_filter[3][3] [2]), .CK(n_53_13), 
      .Q(\buffer[13][3][3] [2]), .QN());
   DFF_X1 \buffer_reg[13][3][3][1]  (.D(\input_filter[3][3] [1]), .CK(n_53_13), 
      .Q(\buffer[13][3][3] [1]), .QN());
   DFF_X1 \buffer_reg[13][3][3][0]  (.D(\input_filter[3][3] [0]), .CK(n_53_13), 
      .Q(\buffer[13][3][3] [0]), .QN());
   DFF_X1 \buffer_reg[14][3][3][15]  (.D(\input_filter[3][3] [15]), .CK(n_53_14), 
      .Q(\buffer[14][3][3] [15]), .QN());
   DFF_X1 \buffer_reg[14][3][3][14]  (.D(\input_filter[3][3] [14]), .CK(n_53_14), 
      .Q(\buffer[14][3][3] [14]), .QN());
   DFF_X1 \buffer_reg[14][3][3][13]  (.D(\input_filter[3][3] [13]), .CK(n_53_14), 
      .Q(\buffer[14][3][3] [13]), .QN());
   DFF_X1 \buffer_reg[14][3][3][12]  (.D(\input_filter[3][3] [12]), .CK(n_53_14), 
      .Q(\buffer[14][3][3] [12]), .QN());
   DFF_X1 \buffer_reg[14][3][3][11]  (.D(\input_filter[3][3] [11]), .CK(n_53_14), 
      .Q(\buffer[14][3][3] [11]), .QN());
   DFF_X1 \buffer_reg[14][3][3][10]  (.D(\input_filter[3][3] [10]), .CK(n_53_14), 
      .Q(\buffer[14][3][3] [10]), .QN());
   DFF_X1 \buffer_reg[14][3][3][9]  (.D(\input_filter[3][3] [9]), .CK(n_53_14), 
      .Q(\buffer[14][3][3] [9]), .QN());
   DFF_X1 \buffer_reg[14][3][3][8]  (.D(\input_filter[3][3] [8]), .CK(n_53_14), 
      .Q(\buffer[14][3][3] [8]), .QN());
   DFF_X1 \buffer_reg[14][3][3][7]  (.D(\input_filter[3][3] [7]), .CK(n_53_14), 
      .Q(\buffer[14][3][3] [7]), .QN());
   DFF_X1 \buffer_reg[14][3][3][6]  (.D(\input_filter[3][3] [6]), .CK(n_53_14), 
      .Q(\buffer[14][3][3] [6]), .QN());
   DFF_X1 \buffer_reg[14][3][3][5]  (.D(\input_filter[3][3] [5]), .CK(n_53_14), 
      .Q(\buffer[14][3][3] [5]), .QN());
   DFF_X1 \buffer_reg[14][3][3][4]  (.D(\input_filter[3][3] [4]), .CK(n_53_14), 
      .Q(\buffer[14][3][3] [4]), .QN());
   DFF_X1 \buffer_reg[14][3][3][3]  (.D(\input_filter[3][3] [3]), .CK(n_53_14), 
      .Q(\buffer[14][3][3] [3]), .QN());
   DFF_X1 \buffer_reg[14][3][3][2]  (.D(\input_filter[3][3] [2]), .CK(n_53_14), 
      .Q(\buffer[14][3][3] [2]), .QN());
   DFF_X1 \buffer_reg[14][3][3][1]  (.D(\input_filter[3][3] [1]), .CK(n_53_14), 
      .Q(\buffer[14][3][3] [1]), .QN());
   DFF_X1 \buffer_reg[14][3][3][0]  (.D(\input_filter[3][3] [0]), .CK(n_53_14), 
      .Q(\buffer[14][3][3] [0]), .QN());
   DFF_X1 \buffer_reg[15][3][3][15]  (.D(\input_filter[3][3] [15]), .CK(n_53_15), 
      .Q(\buffer[15][3][3] [15]), .QN());
   DFF_X1 \buffer_reg[15][3][3][14]  (.D(\input_filter[3][3] [14]), .CK(n_53_15), 
      .Q(\buffer[15][3][3] [14]), .QN());
   DFF_X1 \buffer_reg[15][3][3][13]  (.D(\input_filter[3][3] [13]), .CK(n_53_15), 
      .Q(\buffer[15][3][3] [13]), .QN());
   DFF_X1 \buffer_reg[15][3][3][12]  (.D(\input_filter[3][3] [12]), .CK(n_53_15), 
      .Q(\buffer[15][3][3] [12]), .QN());
   DFF_X1 \buffer_reg[15][3][3][11]  (.D(\input_filter[3][3] [11]), .CK(n_53_15), 
      .Q(\buffer[15][3][3] [11]), .QN());
   DFF_X1 \buffer_reg[15][3][3][10]  (.D(\input_filter[3][3] [10]), .CK(n_53_15), 
      .Q(\buffer[15][3][3] [10]), .QN());
   DFF_X1 \buffer_reg[15][3][3][9]  (.D(\input_filter[3][3] [9]), .CK(n_53_15), 
      .Q(\buffer[15][3][3] [9]), .QN());
   DFF_X1 \buffer_reg[15][3][3][8]  (.D(\input_filter[3][3] [8]), .CK(n_53_15), 
      .Q(\buffer[15][3][3] [8]), .QN());
   DFF_X1 \buffer_reg[15][3][3][7]  (.D(\input_filter[3][3] [7]), .CK(n_53_15), 
      .Q(\buffer[15][3][3] [7]), .QN());
   DFF_X1 \buffer_reg[15][3][3][6]  (.D(\input_filter[3][3] [6]), .CK(n_53_15), 
      .Q(\buffer[15][3][3] [6]), .QN());
   DFF_X1 \buffer_reg[15][3][3][5]  (.D(\input_filter[3][3] [5]), .CK(n_53_15), 
      .Q(\buffer[15][3][3] [5]), .QN());
   DFF_X1 \buffer_reg[15][3][3][4]  (.D(\input_filter[3][3] [4]), .CK(n_53_15), 
      .Q(\buffer[15][3][3] [4]), .QN());
   DFF_X1 \buffer_reg[15][3][3][3]  (.D(\input_filter[3][3] [3]), .CK(n_53_15), 
      .Q(\buffer[15][3][3] [3]), .QN());
   DFF_X1 \buffer_reg[15][3][3][2]  (.D(\input_filter[3][3] [2]), .CK(n_53_15), 
      .Q(\buffer[15][3][3] [2]), .QN());
   DFF_X1 \buffer_reg[15][3][3][1]  (.D(\input_filter[3][3] [1]), .CK(n_53_15), 
      .Q(\buffer[15][3][3] [1]), .QN());
   DFF_X1 \buffer_reg[15][3][3][0]  (.D(\input_filter[3][3] [0]), .CK(n_53_15), 
      .Q(\buffer[15][3][3] [0]), .QN());
   DFF_X1 \buffer_reg[0][3][4][15]  (.D(\input_filter[3][4] [15]), .CK(n_53_0), 
      .Q(\buffer[0][3][4] [15]), .QN());
   DFF_X1 \buffer_reg[0][3][4][14]  (.D(\input_filter[3][4] [14]), .CK(n_53_0), 
      .Q(\buffer[0][3][4] [14]), .QN());
   DFF_X1 \buffer_reg[0][3][4][13]  (.D(\input_filter[3][4] [13]), .CK(n_53_0), 
      .Q(\buffer[0][3][4] [13]), .QN());
   DFF_X1 \buffer_reg[0][3][4][12]  (.D(\input_filter[3][4] [12]), .CK(n_53_0), 
      .Q(\buffer[0][3][4] [12]), .QN());
   DFF_X1 \buffer_reg[0][3][4][11]  (.D(\input_filter[3][4] [11]), .CK(n_53_0), 
      .Q(\buffer[0][3][4] [11]), .QN());
   DFF_X1 \buffer_reg[0][3][4][10]  (.D(\input_filter[3][4] [10]), .CK(n_53_0), 
      .Q(\buffer[0][3][4] [10]), .QN());
   DFF_X1 \buffer_reg[0][3][4][9]  (.D(\input_filter[3][4] [9]), .CK(n_53_0), 
      .Q(\buffer[0][3][4] [9]), .QN());
   DFF_X1 \buffer_reg[0][3][4][8]  (.D(\input_filter[3][4] [8]), .CK(n_53_0), 
      .Q(\buffer[0][3][4] [8]), .QN());
   DFF_X1 \buffer_reg[0][3][4][7]  (.D(\input_filter[3][4] [7]), .CK(n_53_0), 
      .Q(\buffer[0][3][4] [7]), .QN());
   DFF_X1 \buffer_reg[0][3][4][6]  (.D(\input_filter[3][4] [6]), .CK(n_53_0), 
      .Q(\buffer[0][3][4] [6]), .QN());
   DFF_X1 \buffer_reg[0][3][4][5]  (.D(\input_filter[3][4] [5]), .CK(n_53_0), 
      .Q(\buffer[0][3][4] [5]), .QN());
   DFF_X1 \buffer_reg[0][3][4][4]  (.D(\input_filter[3][4] [4]), .CK(n_53_0), 
      .Q(\buffer[0][3][4] [4]), .QN());
   DFF_X1 \buffer_reg[0][3][4][3]  (.D(\input_filter[3][4] [3]), .CK(n_53_0), 
      .Q(\buffer[0][3][4] [3]), .QN());
   DFF_X1 \buffer_reg[0][3][4][2]  (.D(\input_filter[3][4] [2]), .CK(n_53_0), 
      .Q(\buffer[0][3][4] [2]), .QN());
   DFF_X1 \buffer_reg[0][3][4][1]  (.D(\input_filter[3][4] [1]), .CK(n_53_0), 
      .Q(\buffer[0][3][4] [1]), .QN());
   DFF_X1 \buffer_reg[0][3][4][0]  (.D(\input_filter[3][4] [0]), .CK(n_53_0), 
      .Q(\buffer[0][3][4] [0]), .QN());
   DFF_X1 \buffer_reg[1][3][4][15]  (.D(\input_filter[3][4] [15]), .CK(n_53_1), 
      .Q(\buffer[1][3][4] [15]), .QN());
   DFF_X1 \buffer_reg[1][3][4][14]  (.D(\input_filter[3][4] [14]), .CK(n_53_1), 
      .Q(\buffer[1][3][4] [14]), .QN());
   DFF_X1 \buffer_reg[1][3][4][13]  (.D(\input_filter[3][4] [13]), .CK(n_53_1), 
      .Q(\buffer[1][3][4] [13]), .QN());
   DFF_X1 \buffer_reg[1][3][4][12]  (.D(\input_filter[3][4] [12]), .CK(n_53_1), 
      .Q(\buffer[1][3][4] [12]), .QN());
   DFF_X1 \buffer_reg[1][3][4][11]  (.D(\input_filter[3][4] [11]), .CK(n_53_1), 
      .Q(\buffer[1][3][4] [11]), .QN());
   DFF_X1 \buffer_reg[1][3][4][10]  (.D(\input_filter[3][4] [10]), .CK(n_53_1), 
      .Q(\buffer[1][3][4] [10]), .QN());
   DFF_X1 \buffer_reg[1][3][4][9]  (.D(\input_filter[3][4] [9]), .CK(n_53_1), 
      .Q(\buffer[1][3][4] [9]), .QN());
   DFF_X1 \buffer_reg[1][3][4][8]  (.D(\input_filter[3][4] [8]), .CK(n_53_1), 
      .Q(\buffer[1][3][4] [8]), .QN());
   DFF_X1 \buffer_reg[1][3][4][7]  (.D(\input_filter[3][4] [7]), .CK(n_53_1), 
      .Q(\buffer[1][3][4] [7]), .QN());
   DFF_X1 \buffer_reg[1][3][4][6]  (.D(\input_filter[3][4] [6]), .CK(n_53_1), 
      .Q(\buffer[1][3][4] [6]), .QN());
   DFF_X1 \buffer_reg[1][3][4][5]  (.D(\input_filter[3][4] [5]), .CK(n_53_1), 
      .Q(\buffer[1][3][4] [5]), .QN());
   DFF_X1 \buffer_reg[1][3][4][4]  (.D(\input_filter[3][4] [4]), .CK(n_53_1), 
      .Q(\buffer[1][3][4] [4]), .QN());
   DFF_X1 \buffer_reg[1][3][4][3]  (.D(\input_filter[3][4] [3]), .CK(n_53_1), 
      .Q(\buffer[1][3][4] [3]), .QN());
   DFF_X1 \buffer_reg[1][3][4][2]  (.D(\input_filter[3][4] [2]), .CK(n_53_1), 
      .Q(\buffer[1][3][4] [2]), .QN());
   DFF_X1 \buffer_reg[1][3][4][1]  (.D(\input_filter[3][4] [1]), .CK(n_53_1), 
      .Q(\buffer[1][3][4] [1]), .QN());
   DFF_X1 \buffer_reg[1][3][4][0]  (.D(\input_filter[3][4] [0]), .CK(n_53_1), 
      .Q(\buffer[1][3][4] [0]), .QN());
   DFF_X1 \buffer_reg[2][3][4][15]  (.D(\input_filter[3][4] [15]), .CK(n_53_2), 
      .Q(\buffer[2][3][4] [15]), .QN());
   DFF_X1 \buffer_reg[2][3][4][14]  (.D(\input_filter[3][4] [14]), .CK(n_53_2), 
      .Q(\buffer[2][3][4] [14]), .QN());
   DFF_X1 \buffer_reg[2][3][4][13]  (.D(\input_filter[3][4] [13]), .CK(n_53_2), 
      .Q(\buffer[2][3][4] [13]), .QN());
   DFF_X1 \buffer_reg[2][3][4][12]  (.D(\input_filter[3][4] [12]), .CK(n_53_2), 
      .Q(\buffer[2][3][4] [12]), .QN());
   DFF_X1 \buffer_reg[2][3][4][11]  (.D(\input_filter[3][4] [11]), .CK(n_53_2), 
      .Q(\buffer[2][3][4] [11]), .QN());
   DFF_X1 \buffer_reg[2][3][4][10]  (.D(\input_filter[3][4] [10]), .CK(n_53_2), 
      .Q(\buffer[2][3][4] [10]), .QN());
   DFF_X1 \buffer_reg[2][3][4][9]  (.D(\input_filter[3][4] [9]), .CK(n_53_2), 
      .Q(\buffer[2][3][4] [9]), .QN());
   DFF_X1 \buffer_reg[2][3][4][8]  (.D(\input_filter[3][4] [8]), .CK(n_53_2), 
      .Q(\buffer[2][3][4] [8]), .QN());
   DFF_X1 \buffer_reg[2][3][4][7]  (.D(\input_filter[3][4] [7]), .CK(n_53_2), 
      .Q(\buffer[2][3][4] [7]), .QN());
   DFF_X1 \buffer_reg[2][3][4][6]  (.D(\input_filter[3][4] [6]), .CK(n_53_2), 
      .Q(\buffer[2][3][4] [6]), .QN());
   DFF_X1 \buffer_reg[2][3][4][5]  (.D(\input_filter[3][4] [5]), .CK(n_53_2), 
      .Q(\buffer[2][3][4] [5]), .QN());
   DFF_X1 \buffer_reg[2][3][4][4]  (.D(\input_filter[3][4] [4]), .CK(n_53_2), 
      .Q(\buffer[2][3][4] [4]), .QN());
   DFF_X1 \buffer_reg[2][3][4][3]  (.D(\input_filter[3][4] [3]), .CK(n_53_2), 
      .Q(\buffer[2][3][4] [3]), .QN());
   DFF_X1 \buffer_reg[2][3][4][2]  (.D(\input_filter[3][4] [2]), .CK(n_53_2), 
      .Q(\buffer[2][3][4] [2]), .QN());
   DFF_X1 \buffer_reg[2][3][4][1]  (.D(\input_filter[3][4] [1]), .CK(n_53_2), 
      .Q(\buffer[2][3][4] [1]), .QN());
   DFF_X1 \buffer_reg[2][3][4][0]  (.D(\input_filter[3][4] [0]), .CK(n_53_2), 
      .Q(\buffer[2][3][4] [0]), .QN());
   DFF_X1 \buffer_reg[12][4][3][15]  (.D(\input_filter[4][3] [15]), .CK(n_53_12), 
      .Q(\buffer[12][4][3] [15]), .QN());
   DFF_X1 \buffer_reg[12][4][3][14]  (.D(\input_filter[4][3] [14]), .CK(n_53_12), 
      .Q(\buffer[12][4][3] [14]), .QN());
   DFF_X1 \buffer_reg[12][4][3][13]  (.D(\input_filter[4][3] [13]), .CK(n_53_12), 
      .Q(\buffer[12][4][3] [13]), .QN());
   DFF_X1 \buffer_reg[12][4][3][12]  (.D(\input_filter[4][3] [12]), .CK(n_53_12), 
      .Q(\buffer[12][4][3] [12]), .QN());
   DFF_X1 \buffer_reg[12][4][3][11]  (.D(\input_filter[4][3] [11]), .CK(n_53_12), 
      .Q(\buffer[12][4][3] [11]), .QN());
   DFF_X1 \buffer_reg[12][4][3][10]  (.D(\input_filter[4][3] [10]), .CK(n_53_12), 
      .Q(\buffer[12][4][3] [10]), .QN());
   DFF_X1 \buffer_reg[12][4][3][9]  (.D(\input_filter[4][3] [9]), .CK(n_53_12), 
      .Q(\buffer[12][4][3] [9]), .QN());
   DFF_X1 \buffer_reg[12][4][3][8]  (.D(\input_filter[4][3] [8]), .CK(n_53_12), 
      .Q(\buffer[12][4][3] [8]), .QN());
   DFF_X1 \buffer_reg[12][4][3][7]  (.D(\input_filter[4][3] [7]), .CK(n_53_12), 
      .Q(\buffer[12][4][3] [7]), .QN());
   DFF_X1 \buffer_reg[12][4][3][6]  (.D(\input_filter[4][3] [6]), .CK(n_53_12), 
      .Q(\buffer[12][4][3] [6]), .QN());
   DFF_X1 \buffer_reg[12][4][3][5]  (.D(\input_filter[4][3] [5]), .CK(n_53_12), 
      .Q(\buffer[12][4][3] [5]), .QN());
   DFF_X1 \buffer_reg[12][4][3][4]  (.D(\input_filter[4][3] [4]), .CK(n_53_12), 
      .Q(\buffer[12][4][3] [4]), .QN());
   DFF_X1 \buffer_reg[12][4][3][3]  (.D(\input_filter[4][3] [3]), .CK(n_53_12), 
      .Q(\buffer[12][4][3] [3]), .QN());
   DFF_X1 \buffer_reg[12][4][3][2]  (.D(\input_filter[4][3] [2]), .CK(n_53_12), 
      .Q(\buffer[12][4][3] [2]), .QN());
   DFF_X1 \buffer_reg[12][4][3][1]  (.D(\input_filter[4][3] [1]), .CK(n_53_12), 
      .Q(\buffer[12][4][3] [1]), .QN());
   DFF_X1 \buffer_reg[12][4][3][0]  (.D(\input_filter[4][3] [0]), .CK(n_53_12), 
      .Q(\buffer[12][4][3] [0]), .QN());
   DFF_X1 \buffer_reg[11][4][3][15]  (.D(\input_filter[4][3] [15]), .CK(n_53_11), 
      .Q(\buffer[11][4][3] [15]), .QN());
   DFF_X1 \buffer_reg[11][4][3][14]  (.D(\input_filter[4][3] [14]), .CK(n_53_11), 
      .Q(\buffer[11][4][3] [14]), .QN());
   DFF_X1 \buffer_reg[11][4][3][13]  (.D(\input_filter[4][3] [13]), .CK(n_53_11), 
      .Q(\buffer[11][4][3] [13]), .QN());
   DFF_X1 \buffer_reg[11][4][3][12]  (.D(\input_filter[4][3] [12]), .CK(n_53_11), 
      .Q(\buffer[11][4][3] [12]), .QN());
   DFF_X1 \buffer_reg[11][4][3][11]  (.D(\input_filter[4][3] [11]), .CK(n_53_11), 
      .Q(\buffer[11][4][3] [11]), .QN());
   DFF_X1 \buffer_reg[11][4][3][10]  (.D(\input_filter[4][3] [10]), .CK(n_53_11), 
      .Q(\buffer[11][4][3] [10]), .QN());
   DFF_X1 \buffer_reg[11][4][3][9]  (.D(\input_filter[4][3] [9]), .CK(n_53_11), 
      .Q(\buffer[11][4][3] [9]), .QN());
   DFF_X1 \buffer_reg[11][4][3][8]  (.D(\input_filter[4][3] [8]), .CK(n_53_11), 
      .Q(\buffer[11][4][3] [8]), .QN());
   DFF_X1 \buffer_reg[11][4][3][7]  (.D(\input_filter[4][3] [7]), .CK(n_53_11), 
      .Q(\buffer[11][4][3] [7]), .QN());
   DFF_X1 \buffer_reg[11][4][3][6]  (.D(\input_filter[4][3] [6]), .CK(n_53_11), 
      .Q(\buffer[11][4][3] [6]), .QN());
   DFF_X1 \buffer_reg[11][4][3][5]  (.D(\input_filter[4][3] [5]), .CK(n_53_11), 
      .Q(\buffer[11][4][3] [5]), .QN());
   DFF_X1 \buffer_reg[11][4][3][4]  (.D(\input_filter[4][3] [4]), .CK(n_53_11), 
      .Q(\buffer[11][4][3] [4]), .QN());
   DFF_X1 \buffer_reg[11][4][3][3]  (.D(\input_filter[4][3] [3]), .CK(n_53_11), 
      .Q(\buffer[11][4][3] [3]), .QN());
   DFF_X1 \buffer_reg[11][4][3][2]  (.D(\input_filter[4][3] [2]), .CK(n_53_11), 
      .Q(\buffer[11][4][3] [2]), .QN());
   DFF_X1 \buffer_reg[11][4][3][1]  (.D(\input_filter[4][3] [1]), .CK(n_53_11), 
      .Q(\buffer[11][4][3] [1]), .QN());
   DFF_X1 \buffer_reg[11][4][3][0]  (.D(\input_filter[4][3] [0]), .CK(n_53_11), 
      .Q(\buffer[11][4][3] [0]), .QN());
   DFF_X1 \buffer_reg[10][4][3][15]  (.D(\input_filter[4][3] [15]), .CK(n_53_10), 
      .Q(\buffer[10][4][3] [15]), .QN());
   DFF_X1 \buffer_reg[10][4][3][14]  (.D(\input_filter[4][3] [14]), .CK(n_53_10), 
      .Q(\buffer[10][4][3] [14]), .QN());
   DFF_X1 \buffer_reg[10][4][3][13]  (.D(\input_filter[4][3] [13]), .CK(n_53_10), 
      .Q(\buffer[10][4][3] [13]), .QN());
   DFF_X1 \buffer_reg[10][4][3][12]  (.D(\input_filter[4][3] [12]), .CK(n_53_10), 
      .Q(\buffer[10][4][3] [12]), .QN());
   DFF_X1 \buffer_reg[10][4][3][11]  (.D(\input_filter[4][3] [11]), .CK(n_53_10), 
      .Q(\buffer[10][4][3] [11]), .QN());
   DFF_X1 \buffer_reg[10][4][3][10]  (.D(\input_filter[4][3] [10]), .CK(n_53_10), 
      .Q(\buffer[10][4][3] [10]), .QN());
   DFF_X1 \buffer_reg[10][4][3][9]  (.D(\input_filter[4][3] [9]), .CK(n_53_10), 
      .Q(\buffer[10][4][3] [9]), .QN());
   DFF_X1 \buffer_reg[10][4][3][8]  (.D(\input_filter[4][3] [8]), .CK(n_53_10), 
      .Q(\buffer[10][4][3] [8]), .QN());
   DFF_X1 \buffer_reg[10][4][3][7]  (.D(\input_filter[4][3] [7]), .CK(n_53_10), 
      .Q(\buffer[10][4][3] [7]), .QN());
   DFF_X1 \buffer_reg[10][4][3][6]  (.D(\input_filter[4][3] [6]), .CK(n_53_10), 
      .Q(\buffer[10][4][3] [6]), .QN());
   DFF_X1 \buffer_reg[10][4][3][5]  (.D(\input_filter[4][3] [5]), .CK(n_53_10), 
      .Q(\buffer[10][4][3] [5]), .QN());
   DFF_X1 \buffer_reg[10][4][3][4]  (.D(\input_filter[4][3] [4]), .CK(n_53_10), 
      .Q(\buffer[10][4][3] [4]), .QN());
   DFF_X1 \buffer_reg[10][4][3][3]  (.D(\input_filter[4][3] [3]), .CK(n_53_10), 
      .Q(\buffer[10][4][3] [3]), .QN());
   DFF_X1 \buffer_reg[10][4][3][2]  (.D(\input_filter[4][3] [2]), .CK(n_53_10), 
      .Q(\buffer[10][4][3] [2]), .QN());
   DFF_X1 \buffer_reg[10][4][3][1]  (.D(\input_filter[4][3] [1]), .CK(n_53_10), 
      .Q(\buffer[10][4][3] [1]), .QN());
   DFF_X1 \buffer_reg[10][4][3][0]  (.D(\input_filter[4][3] [0]), .CK(n_53_10), 
      .Q(\buffer[10][4][3] [0]), .QN());
   DFF_X1 \buffer_reg[9][4][3][15]  (.D(\input_filter[4][3] [15]), .CK(n_53_9), 
      .Q(\buffer[9][4][3] [15]), .QN());
   DFF_X1 \buffer_reg[9][4][3][14]  (.D(\input_filter[4][3] [14]), .CK(n_53_9), 
      .Q(\buffer[9][4][3] [14]), .QN());
   DFF_X1 \buffer_reg[9][4][3][13]  (.D(\input_filter[4][3] [13]), .CK(n_53_9), 
      .Q(\buffer[9][4][3] [13]), .QN());
   DFF_X1 \buffer_reg[9][4][3][12]  (.D(\input_filter[4][3] [12]), .CK(n_53_9), 
      .Q(\buffer[9][4][3] [12]), .QN());
   DFF_X1 \buffer_reg[9][4][3][11]  (.D(\input_filter[4][3] [11]), .CK(n_53_9), 
      .Q(\buffer[9][4][3] [11]), .QN());
   DFF_X1 \buffer_reg[9][4][3][10]  (.D(\input_filter[4][3] [10]), .CK(n_53_9), 
      .Q(\buffer[9][4][3] [10]), .QN());
   DFF_X1 \buffer_reg[9][4][3][9]  (.D(\input_filter[4][3] [9]), .CK(n_53_9), 
      .Q(\buffer[9][4][3] [9]), .QN());
   DFF_X1 \buffer_reg[9][4][3][8]  (.D(\input_filter[4][3] [8]), .CK(n_53_9), 
      .Q(\buffer[9][4][3] [8]), .QN());
   DFF_X1 \buffer_reg[9][4][3][7]  (.D(\input_filter[4][3] [7]), .CK(n_53_9), 
      .Q(\buffer[9][4][3] [7]), .QN());
   DFF_X1 \buffer_reg[9][4][3][6]  (.D(\input_filter[4][3] [6]), .CK(n_53_9), 
      .Q(\buffer[9][4][3] [6]), .QN());
   DFF_X1 \buffer_reg[9][4][3][5]  (.D(\input_filter[4][3] [5]), .CK(n_53_9), 
      .Q(\buffer[9][4][3] [5]), .QN());
   DFF_X1 \buffer_reg[9][4][3][4]  (.D(\input_filter[4][3] [4]), .CK(n_53_9), 
      .Q(\buffer[9][4][3] [4]), .QN());
   DFF_X1 \buffer_reg[9][4][3][3]  (.D(\input_filter[4][3] [3]), .CK(n_53_9), 
      .Q(\buffer[9][4][3] [3]), .QN());
   DFF_X1 \buffer_reg[9][4][3][2]  (.D(\input_filter[4][3] [2]), .CK(n_53_9), 
      .Q(\buffer[9][4][3] [2]), .QN());
   DFF_X1 \buffer_reg[9][4][3][1]  (.D(\input_filter[4][3] [1]), .CK(n_53_9), 
      .Q(\buffer[9][4][3] [1]), .QN());
   DFF_X1 \buffer_reg[9][4][3][0]  (.D(\input_filter[4][3] [0]), .CK(n_53_9), 
      .Q(\buffer[9][4][3] [0]), .QN());
   DFF_X1 \buffer_reg[8][4][3][15]  (.D(\input_filter[4][3] [15]), .CK(n_53_8), 
      .Q(\buffer[8][4][3] [15]), .QN());
   DFF_X1 \buffer_reg[8][4][3][14]  (.D(\input_filter[4][3] [14]), .CK(n_53_8), 
      .Q(\buffer[8][4][3] [14]), .QN());
   DFF_X1 \buffer_reg[8][4][3][13]  (.D(\input_filter[4][3] [13]), .CK(n_53_8), 
      .Q(\buffer[8][4][3] [13]), .QN());
   DFF_X1 \buffer_reg[8][4][3][12]  (.D(\input_filter[4][3] [12]), .CK(n_53_8), 
      .Q(\buffer[8][4][3] [12]), .QN());
   DFF_X1 \buffer_reg[8][4][3][11]  (.D(\input_filter[4][3] [11]), .CK(n_53_8), 
      .Q(\buffer[8][4][3] [11]), .QN());
   DFF_X1 \buffer_reg[8][4][3][10]  (.D(\input_filter[4][3] [10]), .CK(n_53_8), 
      .Q(\buffer[8][4][3] [10]), .QN());
   DFF_X1 \buffer_reg[8][4][3][9]  (.D(\input_filter[4][3] [9]), .CK(n_53_8), 
      .Q(\buffer[8][4][3] [9]), .QN());
   DFF_X1 \buffer_reg[8][4][3][8]  (.D(\input_filter[4][3] [8]), .CK(n_53_8), 
      .Q(\buffer[8][4][3] [8]), .QN());
   DFF_X1 \buffer_reg[8][4][3][7]  (.D(\input_filter[4][3] [7]), .CK(n_53_8), 
      .Q(\buffer[8][4][3] [7]), .QN());
   DFF_X1 \buffer_reg[8][4][3][6]  (.D(\input_filter[4][3] [6]), .CK(n_53_8), 
      .Q(\buffer[8][4][3] [6]), .QN());
   DFF_X1 \buffer_reg[8][4][3][5]  (.D(\input_filter[4][3] [5]), .CK(n_53_8), 
      .Q(\buffer[8][4][3] [5]), .QN());
   DFF_X1 \buffer_reg[8][4][3][4]  (.D(\input_filter[4][3] [4]), .CK(n_53_8), 
      .Q(\buffer[8][4][3] [4]), .QN());
   DFF_X1 \buffer_reg[8][4][3][3]  (.D(\input_filter[4][3] [3]), .CK(n_53_8), 
      .Q(\buffer[8][4][3] [3]), .QN());
   DFF_X1 \buffer_reg[8][4][3][2]  (.D(\input_filter[4][3] [2]), .CK(n_53_8), 
      .Q(\buffer[8][4][3] [2]), .QN());
   DFF_X1 \buffer_reg[8][4][3][1]  (.D(\input_filter[4][3] [1]), .CK(n_53_8), 
      .Q(\buffer[8][4][3] [1]), .QN());
   DFF_X1 \buffer_reg[8][4][3][0]  (.D(\input_filter[4][3] [0]), .CK(n_53_8), 
      .Q(\buffer[8][4][3] [0]), .QN());
   DFF_X1 \buffer_reg[7][4][3][15]  (.D(\input_filter[4][3] [15]), .CK(n_53_7), 
      .Q(\buffer[7][4][3] [15]), .QN());
   DFF_X1 \buffer_reg[7][4][3][14]  (.D(\input_filter[4][3] [14]), .CK(n_53_7), 
      .Q(\buffer[7][4][3] [14]), .QN());
   DFF_X1 \buffer_reg[7][4][3][13]  (.D(\input_filter[4][3] [13]), .CK(n_53_7), 
      .Q(\buffer[7][4][3] [13]), .QN());
   DFF_X1 \buffer_reg[7][4][3][12]  (.D(\input_filter[4][3] [12]), .CK(n_53_7), 
      .Q(\buffer[7][4][3] [12]), .QN());
   DFF_X1 \buffer_reg[7][4][3][11]  (.D(\input_filter[4][3] [11]), .CK(n_53_7), 
      .Q(\buffer[7][4][3] [11]), .QN());
   DFF_X1 \buffer_reg[7][4][3][10]  (.D(\input_filter[4][3] [10]), .CK(n_53_7), 
      .Q(\buffer[7][4][3] [10]), .QN());
   DFF_X1 \buffer_reg[7][4][3][9]  (.D(\input_filter[4][3] [9]), .CK(n_53_7), 
      .Q(\buffer[7][4][3] [9]), .QN());
   DFF_X1 \buffer_reg[7][4][3][8]  (.D(\input_filter[4][3] [8]), .CK(n_53_7), 
      .Q(\buffer[7][4][3] [8]), .QN());
   DFF_X1 \buffer_reg[7][4][3][7]  (.D(\input_filter[4][3] [7]), .CK(n_53_7), 
      .Q(\buffer[7][4][3] [7]), .QN());
   DFF_X1 \buffer_reg[7][4][3][6]  (.D(\input_filter[4][3] [6]), .CK(n_53_7), 
      .Q(\buffer[7][4][3] [6]), .QN());
   DFF_X1 \buffer_reg[7][4][3][5]  (.D(\input_filter[4][3] [5]), .CK(n_53_7), 
      .Q(\buffer[7][4][3] [5]), .QN());
   DFF_X1 \buffer_reg[7][4][3][4]  (.D(\input_filter[4][3] [4]), .CK(n_53_7), 
      .Q(\buffer[7][4][3] [4]), .QN());
   DFF_X1 \buffer_reg[7][4][3][3]  (.D(\input_filter[4][3] [3]), .CK(n_53_7), 
      .Q(\buffer[7][4][3] [3]), .QN());
   DFF_X1 \buffer_reg[7][4][3][2]  (.D(\input_filter[4][3] [2]), .CK(n_53_7), 
      .Q(\buffer[7][4][3] [2]), .QN());
   DFF_X1 \buffer_reg[7][4][3][1]  (.D(\input_filter[4][3] [1]), .CK(n_53_7), 
      .Q(\buffer[7][4][3] [1]), .QN());
   DFF_X1 \buffer_reg[7][4][3][0]  (.D(\input_filter[4][3] [0]), .CK(n_53_7), 
      .Q(\buffer[7][4][3] [0]), .QN());
   DFF_X1 \buffer_reg[6][4][3][15]  (.D(\input_filter[4][3] [15]), .CK(n_53_6), 
      .Q(\buffer[6][4][3] [15]), .QN());
   DFF_X1 \buffer_reg[6][4][3][14]  (.D(\input_filter[4][3] [14]), .CK(n_53_6), 
      .Q(\buffer[6][4][3] [14]), .QN());
   DFF_X1 \buffer_reg[6][4][3][13]  (.D(\input_filter[4][3] [13]), .CK(n_53_6), 
      .Q(\buffer[6][4][3] [13]), .QN());
   DFF_X1 \buffer_reg[6][4][3][12]  (.D(\input_filter[4][3] [12]), .CK(n_53_6), 
      .Q(\buffer[6][4][3] [12]), .QN());
   DFF_X1 \buffer_reg[6][4][3][11]  (.D(\input_filter[4][3] [11]), .CK(n_53_6), 
      .Q(\buffer[6][4][3] [11]), .QN());
   DFF_X1 \buffer_reg[6][4][3][10]  (.D(\input_filter[4][3] [10]), .CK(n_53_6), 
      .Q(\buffer[6][4][3] [10]), .QN());
   DFF_X1 \buffer_reg[6][4][3][9]  (.D(\input_filter[4][3] [9]), .CK(n_53_6), 
      .Q(\buffer[6][4][3] [9]), .QN());
   DFF_X1 \buffer_reg[6][4][3][8]  (.D(\input_filter[4][3] [8]), .CK(n_53_6), 
      .Q(\buffer[6][4][3] [8]), .QN());
   DFF_X1 \buffer_reg[6][4][3][7]  (.D(\input_filter[4][3] [7]), .CK(n_53_6), 
      .Q(\buffer[6][4][3] [7]), .QN());
   DFF_X1 \buffer_reg[6][4][3][6]  (.D(\input_filter[4][3] [6]), .CK(n_53_6), 
      .Q(\buffer[6][4][3] [6]), .QN());
   DFF_X1 \buffer_reg[6][4][3][5]  (.D(\input_filter[4][3] [5]), .CK(n_53_6), 
      .Q(\buffer[6][4][3] [5]), .QN());
   DFF_X1 \buffer_reg[6][4][3][4]  (.D(\input_filter[4][3] [4]), .CK(n_53_6), 
      .Q(\buffer[6][4][3] [4]), .QN());
   DFF_X1 \buffer_reg[6][4][3][3]  (.D(\input_filter[4][3] [3]), .CK(n_53_6), 
      .Q(\buffer[6][4][3] [3]), .QN());
   DFF_X1 \buffer_reg[6][4][3][2]  (.D(\input_filter[4][3] [2]), .CK(n_53_6), 
      .Q(\buffer[6][4][3] [2]), .QN());
   DFF_X1 \buffer_reg[6][4][3][1]  (.D(\input_filter[4][3] [1]), .CK(n_53_6), 
      .Q(\buffer[6][4][3] [1]), .QN());
   DFF_X1 \buffer_reg[6][4][3][0]  (.D(\input_filter[4][3] [0]), .CK(n_53_6), 
      .Q(\buffer[6][4][3] [0]), .QN());
   DFF_X1 \buffer_reg[5][4][3][15]  (.D(\input_filter[4][3] [15]), .CK(n_53_5), 
      .Q(\buffer[5][4][3] [15]), .QN());
   DFF_X1 \buffer_reg[5][4][3][14]  (.D(\input_filter[4][3] [14]), .CK(n_53_5), 
      .Q(\buffer[5][4][3] [14]), .QN());
   DFF_X1 \buffer_reg[5][4][3][13]  (.D(\input_filter[4][3] [13]), .CK(n_53_5), 
      .Q(\buffer[5][4][3] [13]), .QN());
   DFF_X1 \buffer_reg[5][4][3][12]  (.D(\input_filter[4][3] [12]), .CK(n_53_5), 
      .Q(\buffer[5][4][3] [12]), .QN());
   DFF_X1 \buffer_reg[5][4][3][11]  (.D(\input_filter[4][3] [11]), .CK(n_53_5), 
      .Q(\buffer[5][4][3] [11]), .QN());
   DFF_X1 \buffer_reg[5][4][3][10]  (.D(\input_filter[4][3] [10]), .CK(n_53_5), 
      .Q(\buffer[5][4][3] [10]), .QN());
   DFF_X1 \buffer_reg[5][4][3][9]  (.D(\input_filter[4][3] [9]), .CK(n_53_5), 
      .Q(\buffer[5][4][3] [9]), .QN());
   DFF_X1 \buffer_reg[5][4][3][8]  (.D(\input_filter[4][3] [8]), .CK(n_53_5), 
      .Q(\buffer[5][4][3] [8]), .QN());
   DFF_X1 \buffer_reg[5][4][3][7]  (.D(\input_filter[4][3] [7]), .CK(n_53_5), 
      .Q(\buffer[5][4][3] [7]), .QN());
   DFF_X1 \buffer_reg[5][4][3][6]  (.D(\input_filter[4][3] [6]), .CK(n_53_5), 
      .Q(\buffer[5][4][3] [6]), .QN());
   DFF_X1 \buffer_reg[5][4][3][5]  (.D(\input_filter[4][3] [5]), .CK(n_53_5), 
      .Q(\buffer[5][4][3] [5]), .QN());
   DFF_X1 \buffer_reg[5][4][3][4]  (.D(\input_filter[4][3] [4]), .CK(n_53_5), 
      .Q(\buffer[5][4][3] [4]), .QN());
   DFF_X1 \buffer_reg[5][4][3][3]  (.D(\input_filter[4][3] [3]), .CK(n_53_5), 
      .Q(\buffer[5][4][3] [3]), .QN());
   DFF_X1 \buffer_reg[5][4][3][2]  (.D(\input_filter[4][3] [2]), .CK(n_53_5), 
      .Q(\buffer[5][4][3] [2]), .QN());
   DFF_X1 \buffer_reg[5][4][3][1]  (.D(\input_filter[4][3] [1]), .CK(n_53_5), 
      .Q(\buffer[5][4][3] [1]), .QN());
   DFF_X1 \buffer_reg[5][4][3][0]  (.D(\input_filter[4][3] [0]), .CK(n_53_5), 
      .Q(\buffer[5][4][3] [0]), .QN());
   DFF_X1 \buffer_reg[4][4][3][15]  (.D(\input_filter[4][3] [15]), .CK(n_53_4), 
      .Q(\buffer[4][4][3] [15]), .QN());
   DFF_X1 \buffer_reg[4][4][3][14]  (.D(\input_filter[4][3] [14]), .CK(n_53_4), 
      .Q(\buffer[4][4][3] [14]), .QN());
   DFF_X1 \buffer_reg[4][4][3][13]  (.D(\input_filter[4][3] [13]), .CK(n_53_4), 
      .Q(\buffer[4][4][3] [13]), .QN());
   DFF_X1 \buffer_reg[4][4][3][12]  (.D(\input_filter[4][3] [12]), .CK(n_53_4), 
      .Q(\buffer[4][4][3] [12]), .QN());
   DFF_X1 \buffer_reg[4][4][3][11]  (.D(\input_filter[4][3] [11]), .CK(n_53_4), 
      .Q(\buffer[4][4][3] [11]), .QN());
   DFF_X1 \buffer_reg[4][4][3][10]  (.D(\input_filter[4][3] [10]), .CK(n_53_4), 
      .Q(\buffer[4][4][3] [10]), .QN());
   DFF_X1 \buffer_reg[4][4][3][9]  (.D(\input_filter[4][3] [9]), .CK(n_53_4), 
      .Q(\buffer[4][4][3] [9]), .QN());
   DFF_X1 \buffer_reg[4][4][3][8]  (.D(\input_filter[4][3] [8]), .CK(n_53_4), 
      .Q(\buffer[4][4][3] [8]), .QN());
   DFF_X1 \buffer_reg[4][4][3][7]  (.D(\input_filter[4][3] [7]), .CK(n_53_4), 
      .Q(\buffer[4][4][3] [7]), .QN());
   DFF_X1 \buffer_reg[4][4][3][6]  (.D(\input_filter[4][3] [6]), .CK(n_53_4), 
      .Q(\buffer[4][4][3] [6]), .QN());
   DFF_X1 \buffer_reg[4][4][3][5]  (.D(\input_filter[4][3] [5]), .CK(n_53_4), 
      .Q(\buffer[4][4][3] [5]), .QN());
   DFF_X1 \buffer_reg[4][4][3][4]  (.D(\input_filter[4][3] [4]), .CK(n_53_4), 
      .Q(\buffer[4][4][3] [4]), .QN());
   DFF_X1 \buffer_reg[4][4][3][3]  (.D(\input_filter[4][3] [3]), .CK(n_53_4), 
      .Q(\buffer[4][4][3] [3]), .QN());
   DFF_X1 \buffer_reg[4][4][3][2]  (.D(\input_filter[4][3] [2]), .CK(n_53_4), 
      .Q(\buffer[4][4][3] [2]), .QN());
   DFF_X1 \buffer_reg[4][4][3][1]  (.D(\input_filter[4][3] [1]), .CK(n_53_4), 
      .Q(\buffer[4][4][3] [1]), .QN());
   DFF_X1 \buffer_reg[4][4][3][0]  (.D(\input_filter[4][3] [0]), .CK(n_53_4), 
      .Q(\buffer[4][4][3] [0]), .QN());
   DFF_X1 \buffer_reg[3][3][4][15]  (.D(\input_filter[3][4] [15]), .CK(n_53_3), 
      .Q(\buffer[3][3][4] [15]), .QN());
   DFF_X1 \buffer_reg[3][3][4][14]  (.D(\input_filter[3][4] [14]), .CK(n_53_3), 
      .Q(\buffer[3][3][4] [14]), .QN());
   DFF_X1 \buffer_reg[3][3][4][13]  (.D(\input_filter[3][4] [13]), .CK(n_53_3), 
      .Q(\buffer[3][3][4] [13]), .QN());
   DFF_X1 \buffer_reg[3][3][4][12]  (.D(\input_filter[3][4] [12]), .CK(n_53_3), 
      .Q(\buffer[3][3][4] [12]), .QN());
   DFF_X1 \buffer_reg[3][3][4][11]  (.D(\input_filter[3][4] [11]), .CK(n_53_3), 
      .Q(\buffer[3][3][4] [11]), .QN());
   DFF_X1 \buffer_reg[3][3][4][10]  (.D(\input_filter[3][4] [10]), .CK(n_53_3), 
      .Q(\buffer[3][3][4] [10]), .QN());
   DFF_X1 \buffer_reg[3][3][4][9]  (.D(\input_filter[3][4] [9]), .CK(n_53_3), 
      .Q(\buffer[3][3][4] [9]), .QN());
   DFF_X1 \buffer_reg[3][3][4][8]  (.D(\input_filter[3][4] [8]), .CK(n_53_3), 
      .Q(\buffer[3][3][4] [8]), .QN());
   DFF_X1 \buffer_reg[3][3][4][7]  (.D(\input_filter[3][4] [7]), .CK(n_53_3), 
      .Q(\buffer[3][3][4] [7]), .QN());
   DFF_X1 \buffer_reg[3][3][4][6]  (.D(\input_filter[3][4] [6]), .CK(n_53_3), 
      .Q(\buffer[3][3][4] [6]), .QN());
   DFF_X1 \buffer_reg[3][3][4][5]  (.D(\input_filter[3][4] [5]), .CK(n_53_3), 
      .Q(\buffer[3][3][4] [5]), .QN());
   DFF_X1 \buffer_reg[3][3][4][4]  (.D(\input_filter[3][4] [4]), .CK(n_53_3), 
      .Q(\buffer[3][3][4] [4]), .QN());
   DFF_X1 \buffer_reg[3][3][4][3]  (.D(\input_filter[3][4] [3]), .CK(n_53_3), 
      .Q(\buffer[3][3][4] [3]), .QN());
   DFF_X1 \buffer_reg[3][3][4][2]  (.D(\input_filter[3][4] [2]), .CK(n_53_3), 
      .Q(\buffer[3][3][4] [2]), .QN());
   DFF_X1 \buffer_reg[3][3][4][1]  (.D(\input_filter[3][4] [1]), .CK(n_53_3), 
      .Q(\buffer[3][3][4] [1]), .QN());
   DFF_X1 \buffer_reg[3][3][4][0]  (.D(\input_filter[3][4] [0]), .CK(n_53_3), 
      .Q(\buffer[3][3][4] [0]), .QN());
   DFF_X1 \buffer_reg[4][3][4][15]  (.D(\input_filter[3][4] [15]), .CK(n_53_4), 
      .Q(\buffer[4][3][4] [15]), .QN());
   DFF_X1 \buffer_reg[4][3][4][14]  (.D(\input_filter[3][4] [14]), .CK(n_53_4), 
      .Q(\buffer[4][3][4] [14]), .QN());
   DFF_X1 \buffer_reg[4][3][4][13]  (.D(\input_filter[3][4] [13]), .CK(n_53_4), 
      .Q(\buffer[4][3][4] [13]), .QN());
   DFF_X1 \buffer_reg[4][3][4][12]  (.D(\input_filter[3][4] [12]), .CK(n_53_4), 
      .Q(\buffer[4][3][4] [12]), .QN());
   DFF_X1 \buffer_reg[4][3][4][11]  (.D(\input_filter[3][4] [11]), .CK(n_53_4), 
      .Q(\buffer[4][3][4] [11]), .QN());
   DFF_X1 \buffer_reg[4][3][4][10]  (.D(\input_filter[3][4] [10]), .CK(n_53_4), 
      .Q(\buffer[4][3][4] [10]), .QN());
   DFF_X1 \buffer_reg[4][3][4][9]  (.D(\input_filter[3][4] [9]), .CK(n_53_4), 
      .Q(\buffer[4][3][4] [9]), .QN());
   DFF_X1 \buffer_reg[4][3][4][8]  (.D(\input_filter[3][4] [8]), .CK(n_53_4), 
      .Q(\buffer[4][3][4] [8]), .QN());
   DFF_X1 \buffer_reg[4][3][4][7]  (.D(\input_filter[3][4] [7]), .CK(n_53_4), 
      .Q(\buffer[4][3][4] [7]), .QN());
   DFF_X1 \buffer_reg[4][3][4][6]  (.D(\input_filter[3][4] [6]), .CK(n_53_4), 
      .Q(\buffer[4][3][4] [6]), .QN());
   DFF_X1 \buffer_reg[4][3][4][5]  (.D(\input_filter[3][4] [5]), .CK(n_53_4), 
      .Q(\buffer[4][3][4] [5]), .QN());
   DFF_X1 \buffer_reg[4][3][4][4]  (.D(\input_filter[3][4] [4]), .CK(n_53_4), 
      .Q(\buffer[4][3][4] [4]), .QN());
   DFF_X1 \buffer_reg[4][3][4][3]  (.D(\input_filter[3][4] [3]), .CK(n_53_4), 
      .Q(\buffer[4][3][4] [3]), .QN());
   DFF_X1 \buffer_reg[4][3][4][2]  (.D(\input_filter[3][4] [2]), .CK(n_53_4), 
      .Q(\buffer[4][3][4] [2]), .QN());
   DFF_X1 \buffer_reg[4][3][4][1]  (.D(\input_filter[3][4] [1]), .CK(n_53_4), 
      .Q(\buffer[4][3][4] [1]), .QN());
   DFF_X1 \buffer_reg[4][3][4][0]  (.D(\input_filter[3][4] [0]), .CK(n_53_4), 
      .Q(\buffer[4][3][4] [0]), .QN());
   DFF_X1 \buffer_reg[5][3][4][15]  (.D(\input_filter[3][4] [15]), .CK(n_53_5), 
      .Q(\buffer[5][3][4] [15]), .QN());
   DFF_X1 \buffer_reg[5][3][4][14]  (.D(\input_filter[3][4] [14]), .CK(n_53_5), 
      .Q(\buffer[5][3][4] [14]), .QN());
   DFF_X1 \buffer_reg[5][3][4][13]  (.D(\input_filter[3][4] [13]), .CK(n_53_5), 
      .Q(\buffer[5][3][4] [13]), .QN());
   DFF_X1 \buffer_reg[5][3][4][12]  (.D(\input_filter[3][4] [12]), .CK(n_53_5), 
      .Q(\buffer[5][3][4] [12]), .QN());
   DFF_X1 \buffer_reg[5][3][4][11]  (.D(\input_filter[3][4] [11]), .CK(n_53_5), 
      .Q(\buffer[5][3][4] [11]), .QN());
   DFF_X1 \buffer_reg[5][3][4][10]  (.D(\input_filter[3][4] [10]), .CK(n_53_5), 
      .Q(\buffer[5][3][4] [10]), .QN());
   DFF_X1 \buffer_reg[5][3][4][9]  (.D(\input_filter[3][4] [9]), .CK(n_53_5), 
      .Q(\buffer[5][3][4] [9]), .QN());
   DFF_X1 \buffer_reg[5][3][4][8]  (.D(\input_filter[3][4] [8]), .CK(n_53_5), 
      .Q(\buffer[5][3][4] [8]), .QN());
   DFF_X1 \buffer_reg[5][3][4][7]  (.D(\input_filter[3][4] [7]), .CK(n_53_5), 
      .Q(\buffer[5][3][4] [7]), .QN());
   DFF_X1 \buffer_reg[5][3][4][6]  (.D(\input_filter[3][4] [6]), .CK(n_53_5), 
      .Q(\buffer[5][3][4] [6]), .QN());
   DFF_X1 \buffer_reg[5][3][4][5]  (.D(\input_filter[3][4] [5]), .CK(n_53_5), 
      .Q(\buffer[5][3][4] [5]), .QN());
   DFF_X1 \buffer_reg[5][3][4][4]  (.D(\input_filter[3][4] [4]), .CK(n_53_5), 
      .Q(\buffer[5][3][4] [4]), .QN());
   DFF_X1 \buffer_reg[5][3][4][3]  (.D(\input_filter[3][4] [3]), .CK(n_53_5), 
      .Q(\buffer[5][3][4] [3]), .QN());
   DFF_X1 \buffer_reg[5][3][4][2]  (.D(\input_filter[3][4] [2]), .CK(n_53_5), 
      .Q(\buffer[5][3][4] [2]), .QN());
   DFF_X1 \buffer_reg[5][3][4][1]  (.D(\input_filter[3][4] [1]), .CK(n_53_5), 
      .Q(\buffer[5][3][4] [1]), .QN());
   DFF_X1 \buffer_reg[5][3][4][0]  (.D(\input_filter[3][4] [0]), .CK(n_53_5), 
      .Q(\buffer[5][3][4] [0]), .QN());
   DFF_X1 \buffer_reg[0][4][3][15]  (.D(\input_filter[4][3] [15]), .CK(n_53_0), 
      .Q(\buffer[0][4][3] [15]), .QN());
   DFF_X1 \buffer_reg[0][4][3][14]  (.D(\input_filter[4][3] [14]), .CK(n_53_0), 
      .Q(\buffer[0][4][3] [14]), .QN());
   DFF_X1 \buffer_reg[0][4][3][13]  (.D(\input_filter[4][3] [13]), .CK(n_53_0), 
      .Q(\buffer[0][4][3] [13]), .QN());
   DFF_X1 \buffer_reg[0][4][3][12]  (.D(\input_filter[4][3] [12]), .CK(n_53_0), 
      .Q(\buffer[0][4][3] [12]), .QN());
   DFF_X1 \buffer_reg[0][4][3][11]  (.D(\input_filter[4][3] [11]), .CK(n_53_0), 
      .Q(\buffer[0][4][3] [11]), .QN());
   DFF_X1 \buffer_reg[0][4][3][10]  (.D(\input_filter[4][3] [10]), .CK(n_53_0), 
      .Q(\buffer[0][4][3] [10]), .QN());
   DFF_X1 \buffer_reg[0][4][3][9]  (.D(\input_filter[4][3] [9]), .CK(n_53_0), 
      .Q(\buffer[0][4][3] [9]), .QN());
   DFF_X1 \buffer_reg[0][4][3][8]  (.D(\input_filter[4][3] [8]), .CK(n_53_0), 
      .Q(\buffer[0][4][3] [8]), .QN());
   DFF_X1 \buffer_reg[0][4][3][7]  (.D(\input_filter[4][3] [7]), .CK(n_53_0), 
      .Q(\buffer[0][4][3] [7]), .QN());
   DFF_X1 \buffer_reg[0][4][3][6]  (.D(\input_filter[4][3] [6]), .CK(n_53_0), 
      .Q(\buffer[0][4][3] [6]), .QN());
   DFF_X1 \buffer_reg[0][4][3][5]  (.D(\input_filter[4][3] [5]), .CK(n_53_0), 
      .Q(\buffer[0][4][3] [5]), .QN());
   DFF_X1 \buffer_reg[0][4][3][4]  (.D(\input_filter[4][3] [4]), .CK(n_53_0), 
      .Q(\buffer[0][4][3] [4]), .QN());
   DFF_X1 \buffer_reg[0][4][3][3]  (.D(\input_filter[4][3] [3]), .CK(n_53_0), 
      .Q(\buffer[0][4][3] [3]), .QN());
   DFF_X1 \buffer_reg[0][4][3][2]  (.D(\input_filter[4][3] [2]), .CK(n_53_0), 
      .Q(\buffer[0][4][3] [2]), .QN());
   DFF_X1 \buffer_reg[0][4][3][1]  (.D(\input_filter[4][3] [1]), .CK(n_53_0), 
      .Q(\buffer[0][4][3] [1]), .QN());
   DFF_X1 \buffer_reg[0][4][3][0]  (.D(\input_filter[4][3] [0]), .CK(n_53_0), 
      .Q(\buffer[0][4][3] [0]), .QN());
   DFF_X1 \buffer_reg[15][4][2][15]  (.D(\input_filter[4][2] [15]), .CK(n_53_15), 
      .Q(\buffer[15][4][2] [15]), .QN());
   DFF_X1 \buffer_reg[15][4][2][14]  (.D(\input_filter[4][2] [14]), .CK(n_53_15), 
      .Q(\buffer[15][4][2] [14]), .QN());
   DFF_X1 \buffer_reg[15][4][2][13]  (.D(\input_filter[4][2] [13]), .CK(n_53_15), 
      .Q(\buffer[15][4][2] [13]), .QN());
   DFF_X1 \buffer_reg[15][4][2][12]  (.D(\input_filter[4][2] [12]), .CK(n_53_15), 
      .Q(\buffer[15][4][2] [12]), .QN());
   DFF_X1 \buffer_reg[15][4][2][11]  (.D(\input_filter[4][2] [11]), .CK(n_53_15), 
      .Q(\buffer[15][4][2] [11]), .QN());
   DFF_X1 \buffer_reg[15][4][2][10]  (.D(\input_filter[4][2] [10]), .CK(n_53_15), 
      .Q(\buffer[15][4][2] [10]), .QN());
   DFF_X1 \buffer_reg[15][4][2][9]  (.D(\input_filter[4][2] [9]), .CK(n_53_15), 
      .Q(\buffer[15][4][2] [9]), .QN());
   DFF_X1 \buffer_reg[15][4][2][8]  (.D(\input_filter[4][2] [8]), .CK(n_53_15), 
      .Q(\buffer[15][4][2] [8]), .QN());
   DFF_X1 \buffer_reg[15][4][2][7]  (.D(\input_filter[4][2] [7]), .CK(n_53_15), 
      .Q(\buffer[15][4][2] [7]), .QN());
   DFF_X1 \buffer_reg[15][4][2][6]  (.D(\input_filter[4][2] [6]), .CK(n_53_15), 
      .Q(\buffer[15][4][2] [6]), .QN());
   DFF_X1 \buffer_reg[15][4][2][5]  (.D(\input_filter[4][2] [5]), .CK(n_53_15), 
      .Q(\buffer[15][4][2] [5]), .QN());
   DFF_X1 \buffer_reg[15][4][2][4]  (.D(\input_filter[4][2] [4]), .CK(n_53_15), 
      .Q(\buffer[15][4][2] [4]), .QN());
   DFF_X1 \buffer_reg[15][4][2][3]  (.D(\input_filter[4][2] [3]), .CK(n_53_15), 
      .Q(\buffer[15][4][2] [3]), .QN());
   DFF_X1 \buffer_reg[15][4][2][2]  (.D(\input_filter[4][2] [2]), .CK(n_53_15), 
      .Q(\buffer[15][4][2] [2]), .QN());
   DFF_X1 \buffer_reg[15][4][2][1]  (.D(\input_filter[4][2] [1]), .CK(n_53_15), 
      .Q(\buffer[15][4][2] [1]), .QN());
   DFF_X1 \buffer_reg[15][4][2][0]  (.D(\input_filter[4][2] [0]), .CK(n_53_15), 
      .Q(\buffer[15][4][2] [0]), .QN());
   DFF_X1 \buffer_reg[14][4][2][15]  (.D(\input_filter[4][2] [15]), .CK(n_53_14), 
      .Q(\buffer[14][4][2] [15]), .QN());
   DFF_X1 \buffer_reg[14][4][2][14]  (.D(\input_filter[4][2] [14]), .CK(n_53_14), 
      .Q(\buffer[14][4][2] [14]), .QN());
   DFF_X1 \buffer_reg[14][4][2][13]  (.D(\input_filter[4][2] [13]), .CK(n_53_14), 
      .Q(\buffer[14][4][2] [13]), .QN());
   DFF_X1 \buffer_reg[14][4][2][12]  (.D(\input_filter[4][2] [12]), .CK(n_53_14), 
      .Q(\buffer[14][4][2] [12]), .QN());
   DFF_X1 \buffer_reg[14][4][2][11]  (.D(\input_filter[4][2] [11]), .CK(n_53_14), 
      .Q(\buffer[14][4][2] [11]), .QN());
   DFF_X1 \buffer_reg[14][4][2][10]  (.D(\input_filter[4][2] [10]), .CK(n_53_14), 
      .Q(\buffer[14][4][2] [10]), .QN());
   DFF_X1 \buffer_reg[14][4][2][9]  (.D(\input_filter[4][2] [9]), .CK(n_53_14), 
      .Q(\buffer[14][4][2] [9]), .QN());
   DFF_X1 \buffer_reg[14][4][2][8]  (.D(\input_filter[4][2] [8]), .CK(n_53_14), 
      .Q(\buffer[14][4][2] [8]), .QN());
   DFF_X1 \buffer_reg[14][4][2][7]  (.D(\input_filter[4][2] [7]), .CK(n_53_14), 
      .Q(\buffer[14][4][2] [7]), .QN());
   DFF_X1 \buffer_reg[14][4][2][6]  (.D(\input_filter[4][2] [6]), .CK(n_53_14), 
      .Q(\buffer[14][4][2] [6]), .QN());
   DFF_X1 \buffer_reg[14][4][2][5]  (.D(\input_filter[4][2] [5]), .CK(n_53_14), 
      .Q(\buffer[14][4][2] [5]), .QN());
   DFF_X1 \buffer_reg[14][4][2][4]  (.D(\input_filter[4][2] [4]), .CK(n_53_14), 
      .Q(\buffer[14][4][2] [4]), .QN());
   DFF_X1 \buffer_reg[14][4][2][3]  (.D(\input_filter[4][2] [3]), .CK(n_53_14), 
      .Q(\buffer[14][4][2] [3]), .QN());
   DFF_X1 \buffer_reg[14][4][2][2]  (.D(\input_filter[4][2] [2]), .CK(n_53_14), 
      .Q(\buffer[14][4][2] [2]), .QN());
   DFF_X1 \buffer_reg[14][4][2][1]  (.D(\input_filter[4][2] [1]), .CK(n_53_14), 
      .Q(\buffer[14][4][2] [1]), .QN());
   DFF_X1 \buffer_reg[14][4][2][0]  (.D(\input_filter[4][2] [0]), .CK(n_53_14), 
      .Q(\buffer[14][4][2] [0]), .QN());
   DFF_X1 \buffer_reg[13][4][2][15]  (.D(\input_filter[4][2] [15]), .CK(n_53_13), 
      .Q(\buffer[13][4][2] [15]), .QN());
   DFF_X1 \buffer_reg[13][4][2][14]  (.D(\input_filter[4][2] [14]), .CK(n_53_13), 
      .Q(\buffer[13][4][2] [14]), .QN());
   DFF_X1 \buffer_reg[13][4][2][13]  (.D(\input_filter[4][2] [13]), .CK(n_53_13), 
      .Q(\buffer[13][4][2] [13]), .QN());
   DFF_X1 \buffer_reg[13][4][2][12]  (.D(\input_filter[4][2] [12]), .CK(n_53_13), 
      .Q(\buffer[13][4][2] [12]), .QN());
   DFF_X1 \buffer_reg[13][4][2][11]  (.D(\input_filter[4][2] [11]), .CK(n_53_13), 
      .Q(\buffer[13][4][2] [11]), .QN());
   DFF_X1 \buffer_reg[13][4][2][10]  (.D(\input_filter[4][2] [10]), .CK(n_53_13), 
      .Q(\buffer[13][4][2] [10]), .QN());
   DFF_X1 \buffer_reg[13][4][2][9]  (.D(\input_filter[4][2] [9]), .CK(n_53_13), 
      .Q(\buffer[13][4][2] [9]), .QN());
   DFF_X1 \buffer_reg[13][4][2][8]  (.D(\input_filter[4][2] [8]), .CK(n_53_13), 
      .Q(\buffer[13][4][2] [8]), .QN());
   DFF_X1 \buffer_reg[13][4][2][7]  (.D(\input_filter[4][2] [7]), .CK(n_53_13), 
      .Q(\buffer[13][4][2] [7]), .QN());
   DFF_X1 \buffer_reg[13][4][2][6]  (.D(\input_filter[4][2] [6]), .CK(n_53_13), 
      .Q(\buffer[13][4][2] [6]), .QN());
   DFF_X1 \buffer_reg[13][4][2][5]  (.D(\input_filter[4][2] [5]), .CK(n_53_13), 
      .Q(\buffer[13][4][2] [5]), .QN());
   DFF_X1 \buffer_reg[13][4][2][4]  (.D(\input_filter[4][2] [4]), .CK(n_53_13), 
      .Q(\buffer[13][4][2] [4]), .QN());
   DFF_X1 \buffer_reg[13][4][2][3]  (.D(\input_filter[4][2] [3]), .CK(n_53_13), 
      .Q(\buffer[13][4][2] [3]), .QN());
   DFF_X1 \buffer_reg[13][4][2][2]  (.D(\input_filter[4][2] [2]), .CK(n_53_13), 
      .Q(\buffer[13][4][2] [2]), .QN());
   DFF_X1 \buffer_reg[13][4][2][1]  (.D(\input_filter[4][2] [1]), .CK(n_53_13), 
      .Q(\buffer[13][4][2] [1]), .QN());
   DFF_X1 \buffer_reg[13][4][2][0]  (.D(\input_filter[4][2] [0]), .CK(n_53_13), 
      .Q(\buffer[13][4][2] [0]), .QN());
   DFF_X1 \buffer_reg[12][4][2][15]  (.D(\input_filter[4][2] [15]), .CK(n_53_12), 
      .Q(\buffer[12][4][2] [15]), .QN());
   DFF_X1 \buffer_reg[12][4][2][14]  (.D(\input_filter[4][2] [14]), .CK(n_53_12), 
      .Q(\buffer[12][4][2] [14]), .QN());
   DFF_X1 \buffer_reg[12][4][2][13]  (.D(\input_filter[4][2] [13]), .CK(n_53_12), 
      .Q(\buffer[12][4][2] [13]), .QN());
   DFF_X1 \buffer_reg[12][4][2][12]  (.D(\input_filter[4][2] [12]), .CK(n_53_12), 
      .Q(\buffer[12][4][2] [12]), .QN());
   DFF_X1 \buffer_reg[12][4][2][11]  (.D(\input_filter[4][2] [11]), .CK(n_53_12), 
      .Q(\buffer[12][4][2] [11]), .QN());
   DFF_X1 \buffer_reg[12][4][2][10]  (.D(\input_filter[4][2] [10]), .CK(n_53_12), 
      .Q(\buffer[12][4][2] [10]), .QN());
   DFF_X1 \buffer_reg[12][4][2][9]  (.D(\input_filter[4][2] [9]), .CK(n_53_12), 
      .Q(\buffer[12][4][2] [9]), .QN());
   DFF_X1 \buffer_reg[12][4][2][8]  (.D(\input_filter[4][2] [8]), .CK(n_53_12), 
      .Q(\buffer[12][4][2] [8]), .QN());
   DFF_X1 \buffer_reg[12][4][2][7]  (.D(\input_filter[4][2] [7]), .CK(n_53_12), 
      .Q(\buffer[12][4][2] [7]), .QN());
   DFF_X1 \buffer_reg[12][4][2][6]  (.D(\input_filter[4][2] [6]), .CK(n_53_12), 
      .Q(\buffer[12][4][2] [6]), .QN());
   DFF_X1 \buffer_reg[12][4][2][5]  (.D(\input_filter[4][2] [5]), .CK(n_53_12), 
      .Q(\buffer[12][4][2] [5]), .QN());
   DFF_X1 \buffer_reg[12][4][2][4]  (.D(\input_filter[4][2] [4]), .CK(n_53_12), 
      .Q(\buffer[12][4][2] [4]), .QN());
   DFF_X1 \buffer_reg[12][4][2][3]  (.D(\input_filter[4][2] [3]), .CK(n_53_12), 
      .Q(\buffer[12][4][2] [3]), .QN());
   DFF_X1 \buffer_reg[12][4][2][2]  (.D(\input_filter[4][2] [2]), .CK(n_53_12), 
      .Q(\buffer[12][4][2] [2]), .QN());
   DFF_X1 \buffer_reg[12][4][2][1]  (.D(\input_filter[4][2] [1]), .CK(n_53_12), 
      .Q(\buffer[12][4][2] [1]), .QN());
   DFF_X1 \buffer_reg[12][4][2][0]  (.D(\input_filter[4][2] [0]), .CK(n_53_12), 
      .Q(\buffer[12][4][2] [0]), .QN());
   DFF_X1 \buffer_reg[11][4][2][15]  (.D(\input_filter[4][2] [15]), .CK(n_53_11), 
      .Q(\buffer[11][4][2] [15]), .QN());
   DFF_X1 \buffer_reg[11][4][2][14]  (.D(\input_filter[4][2] [14]), .CK(n_53_11), 
      .Q(\buffer[11][4][2] [14]), .QN());
   DFF_X1 \buffer_reg[11][4][2][13]  (.D(\input_filter[4][2] [13]), .CK(n_53_11), 
      .Q(\buffer[11][4][2] [13]), .QN());
   DFF_X1 \buffer_reg[11][4][2][12]  (.D(\input_filter[4][2] [12]), .CK(n_53_11), 
      .Q(\buffer[11][4][2] [12]), .QN());
   DFF_X1 \buffer_reg[11][4][2][11]  (.D(\input_filter[4][2] [11]), .CK(n_53_11), 
      .Q(\buffer[11][4][2] [11]), .QN());
   DFF_X1 \buffer_reg[11][4][2][10]  (.D(\input_filter[4][2] [10]), .CK(n_53_11), 
      .Q(\buffer[11][4][2] [10]), .QN());
   DFF_X1 \buffer_reg[11][4][2][9]  (.D(\input_filter[4][2] [9]), .CK(n_53_11), 
      .Q(\buffer[11][4][2] [9]), .QN());
   DFF_X1 \buffer_reg[11][4][2][8]  (.D(\input_filter[4][2] [8]), .CK(n_53_11), 
      .Q(\buffer[11][4][2] [8]), .QN());
   DFF_X1 \buffer_reg[11][4][2][7]  (.D(\input_filter[4][2] [7]), .CK(n_53_11), 
      .Q(\buffer[11][4][2] [7]), .QN());
   DFF_X1 \buffer_reg[11][4][2][6]  (.D(\input_filter[4][2] [6]), .CK(n_53_11), 
      .Q(\buffer[11][4][2] [6]), .QN());
   DFF_X1 \buffer_reg[11][4][2][5]  (.D(\input_filter[4][2] [5]), .CK(n_53_11), 
      .Q(\buffer[11][4][2] [5]), .QN());
   DFF_X1 \buffer_reg[11][4][2][4]  (.D(\input_filter[4][2] [4]), .CK(n_53_11), 
      .Q(\buffer[11][4][2] [4]), .QN());
   DFF_X1 \buffer_reg[11][4][2][3]  (.D(\input_filter[4][2] [3]), .CK(n_53_11), 
      .Q(\buffer[11][4][2] [3]), .QN());
   DFF_X1 \buffer_reg[11][4][2][2]  (.D(\input_filter[4][2] [2]), .CK(n_53_11), 
      .Q(\buffer[11][4][2] [2]), .QN());
   DFF_X1 \buffer_reg[11][4][2][1]  (.D(\input_filter[4][2] [1]), .CK(n_53_11), 
      .Q(\buffer[11][4][2] [1]), .QN());
   DFF_X1 \buffer_reg[11][4][2][0]  (.D(\input_filter[4][2] [0]), .CK(n_53_11), 
      .Q(\buffer[11][4][2] [0]), .QN());
   DFF_X1 \buffer_reg[10][4][2][15]  (.D(\input_filter[4][2] [15]), .CK(n_53_10), 
      .Q(\buffer[10][4][2] [15]), .QN());
   DFF_X1 \buffer_reg[10][4][2][14]  (.D(\input_filter[4][2] [14]), .CK(n_53_10), 
      .Q(\buffer[10][4][2] [14]), .QN());
   DFF_X1 \buffer_reg[10][4][2][13]  (.D(\input_filter[4][2] [13]), .CK(n_53_10), 
      .Q(\buffer[10][4][2] [13]), .QN());
   DFF_X1 \buffer_reg[10][4][2][12]  (.D(\input_filter[4][2] [12]), .CK(n_53_10), 
      .Q(\buffer[10][4][2] [12]), .QN());
   DFF_X1 \buffer_reg[10][4][2][11]  (.D(\input_filter[4][2] [11]), .CK(n_53_10), 
      .Q(\buffer[10][4][2] [11]), .QN());
   DFF_X1 \buffer_reg[10][4][2][10]  (.D(\input_filter[4][2] [10]), .CK(n_53_10), 
      .Q(\buffer[10][4][2] [10]), .QN());
   DFF_X1 \buffer_reg[10][4][2][9]  (.D(\input_filter[4][2] [9]), .CK(n_53_10), 
      .Q(\buffer[10][4][2] [9]), .QN());
   DFF_X1 \buffer_reg[10][4][2][8]  (.D(\input_filter[4][2] [8]), .CK(n_53_10), 
      .Q(\buffer[10][4][2] [8]), .QN());
   DFF_X1 \buffer_reg[10][4][2][7]  (.D(\input_filter[4][2] [7]), .CK(n_53_10), 
      .Q(\buffer[10][4][2] [7]), .QN());
   DFF_X1 \buffer_reg[10][4][2][6]  (.D(\input_filter[4][2] [6]), .CK(n_53_10), 
      .Q(\buffer[10][4][2] [6]), .QN());
   DFF_X1 \buffer_reg[10][4][2][5]  (.D(\input_filter[4][2] [5]), .CK(n_53_10), 
      .Q(\buffer[10][4][2] [5]), .QN());
   DFF_X1 \buffer_reg[10][4][2][4]  (.D(\input_filter[4][2] [4]), .CK(n_53_10), 
      .Q(\buffer[10][4][2] [4]), .QN());
   DFF_X1 \buffer_reg[10][4][2][3]  (.D(\input_filter[4][2] [3]), .CK(n_53_10), 
      .Q(\buffer[10][4][2] [3]), .QN());
   DFF_X1 \buffer_reg[10][4][2][2]  (.D(\input_filter[4][2] [2]), .CK(n_53_10), 
      .Q(\buffer[10][4][2] [2]), .QN());
   DFF_X1 \buffer_reg[10][4][2][1]  (.D(\input_filter[4][2] [1]), .CK(n_53_10), 
      .Q(\buffer[10][4][2] [1]), .QN());
   DFF_X1 \buffer_reg[10][4][2][0]  (.D(\input_filter[4][2] [0]), .CK(n_53_10), 
      .Q(\buffer[10][4][2] [0]), .QN());
   DFF_X1 \buffer_reg[9][4][2][15]  (.D(\input_filter[4][2] [15]), .CK(n_53_9), 
      .Q(\buffer[9][4][2] [15]), .QN());
   DFF_X1 \buffer_reg[9][4][2][14]  (.D(\input_filter[4][2] [14]), .CK(n_53_9), 
      .Q(\buffer[9][4][2] [14]), .QN());
   DFF_X1 \buffer_reg[9][4][2][13]  (.D(\input_filter[4][2] [13]), .CK(n_53_9), 
      .Q(\buffer[9][4][2] [13]), .QN());
   DFF_X1 \buffer_reg[9][4][2][12]  (.D(\input_filter[4][2] [12]), .CK(n_53_9), 
      .Q(\buffer[9][4][2] [12]), .QN());
   DFF_X1 \buffer_reg[9][4][2][11]  (.D(\input_filter[4][2] [11]), .CK(n_53_9), 
      .Q(\buffer[9][4][2] [11]), .QN());
   DFF_X1 \buffer_reg[9][4][2][10]  (.D(\input_filter[4][2] [10]), .CK(n_53_9), 
      .Q(\buffer[9][4][2] [10]), .QN());
   DFF_X1 \buffer_reg[9][4][2][9]  (.D(\input_filter[4][2] [9]), .CK(n_53_9), 
      .Q(\buffer[9][4][2] [9]), .QN());
   DFF_X1 \buffer_reg[9][4][2][8]  (.D(\input_filter[4][2] [8]), .CK(n_53_9), 
      .Q(\buffer[9][4][2] [8]), .QN());
   DFF_X1 \buffer_reg[9][4][2][7]  (.D(\input_filter[4][2] [7]), .CK(n_53_9), 
      .Q(\buffer[9][4][2] [7]), .QN());
   DFF_X1 \buffer_reg[9][4][2][6]  (.D(\input_filter[4][2] [6]), .CK(n_53_9), 
      .Q(\buffer[9][4][2] [6]), .QN());
   DFF_X1 \buffer_reg[9][4][2][5]  (.D(\input_filter[4][2] [5]), .CK(n_53_9), 
      .Q(\buffer[9][4][2] [5]), .QN());
   DFF_X1 \buffer_reg[9][4][2][4]  (.D(\input_filter[4][2] [4]), .CK(n_53_9), 
      .Q(\buffer[9][4][2] [4]), .QN());
   DFF_X1 \buffer_reg[9][4][2][3]  (.D(\input_filter[4][2] [3]), .CK(n_53_9), 
      .Q(\buffer[9][4][2] [3]), .QN());
   DFF_X1 \buffer_reg[9][4][2][2]  (.D(\input_filter[4][2] [2]), .CK(n_53_9), 
      .Q(\buffer[9][4][2] [2]), .QN());
   DFF_X1 \buffer_reg[9][4][2][1]  (.D(\input_filter[4][2] [1]), .CK(n_53_9), 
      .Q(\buffer[9][4][2] [1]), .QN());
   DFF_X1 \buffer_reg[9][4][2][0]  (.D(\input_filter[4][2] [0]), .CK(n_53_9), 
      .Q(\buffer[9][4][2] [0]), .QN());
   DFF_X1 \buffer_reg[8][4][2][15]  (.D(\input_filter[4][2] [15]), .CK(n_53_8), 
      .Q(\buffer[8][4][2] [15]), .QN());
   DFF_X1 \buffer_reg[8][4][2][14]  (.D(\input_filter[4][2] [14]), .CK(n_53_8), 
      .Q(\buffer[8][4][2] [14]), .QN());
   DFF_X1 \buffer_reg[8][4][2][13]  (.D(\input_filter[4][2] [13]), .CK(n_53_8), 
      .Q(\buffer[8][4][2] [13]), .QN());
   DFF_X1 \buffer_reg[8][4][2][12]  (.D(\input_filter[4][2] [12]), .CK(n_53_8), 
      .Q(\buffer[8][4][2] [12]), .QN());
   DFF_X1 \buffer_reg[8][4][2][11]  (.D(\input_filter[4][2] [11]), .CK(n_53_8), 
      .Q(\buffer[8][4][2] [11]), .QN());
   DFF_X1 \buffer_reg[8][4][2][10]  (.D(\input_filter[4][2] [10]), .CK(n_53_8), 
      .Q(\buffer[8][4][2] [10]), .QN());
   DFF_X1 \buffer_reg[8][4][2][9]  (.D(\input_filter[4][2] [9]), .CK(n_53_8), 
      .Q(\buffer[8][4][2] [9]), .QN());
   DFF_X1 \buffer_reg[8][4][2][8]  (.D(\input_filter[4][2] [8]), .CK(n_53_8), 
      .Q(\buffer[8][4][2] [8]), .QN());
   DFF_X1 \buffer_reg[8][4][2][7]  (.D(\input_filter[4][2] [7]), .CK(n_53_8), 
      .Q(\buffer[8][4][2] [7]), .QN());
   DFF_X1 \buffer_reg[8][4][2][6]  (.D(\input_filter[4][2] [6]), .CK(n_53_8), 
      .Q(\buffer[8][4][2] [6]), .QN());
   DFF_X1 \buffer_reg[8][4][2][5]  (.D(\input_filter[4][2] [5]), .CK(n_53_8), 
      .Q(\buffer[8][4][2] [5]), .QN());
   DFF_X1 \buffer_reg[8][4][2][4]  (.D(\input_filter[4][2] [4]), .CK(n_53_8), 
      .Q(\buffer[8][4][2] [4]), .QN());
   DFF_X1 \buffer_reg[8][4][2][3]  (.D(\input_filter[4][2] [3]), .CK(n_53_8), 
      .Q(\buffer[8][4][2] [3]), .QN());
   DFF_X1 \buffer_reg[8][4][2][2]  (.D(\input_filter[4][2] [2]), .CK(n_53_8), 
      .Q(\buffer[8][4][2] [2]), .QN());
   DFF_X1 \buffer_reg[8][4][2][1]  (.D(\input_filter[4][2] [1]), .CK(n_53_8), 
      .Q(\buffer[8][4][2] [1]), .QN());
   DFF_X1 \buffer_reg[8][4][2][0]  (.D(\input_filter[4][2] [0]), .CK(n_53_8), 
      .Q(\buffer[8][4][2] [0]), .QN());
   DFF_X1 \buffer_reg[7][4][2][15]  (.D(\input_filter[4][2] [15]), .CK(n_53_7), 
      .Q(\buffer[7][4][2] [15]), .QN());
   DFF_X1 \buffer_reg[7][4][2][14]  (.D(\input_filter[4][2] [14]), .CK(n_53_7), 
      .Q(\buffer[7][4][2] [14]), .QN());
   DFF_X1 \buffer_reg[7][4][2][13]  (.D(\input_filter[4][2] [13]), .CK(n_53_7), 
      .Q(\buffer[7][4][2] [13]), .QN());
   DFF_X1 \buffer_reg[7][4][2][12]  (.D(\input_filter[4][2] [12]), .CK(n_53_7), 
      .Q(\buffer[7][4][2] [12]), .QN());
   DFF_X1 \buffer_reg[7][4][2][11]  (.D(\input_filter[4][2] [11]), .CK(n_53_7), 
      .Q(\buffer[7][4][2] [11]), .QN());
   DFF_X1 \buffer_reg[7][4][2][10]  (.D(\input_filter[4][2] [10]), .CK(n_53_7), 
      .Q(\buffer[7][4][2] [10]), .QN());
   DFF_X1 \buffer_reg[7][4][2][9]  (.D(\input_filter[4][2] [9]), .CK(n_53_7), 
      .Q(\buffer[7][4][2] [9]), .QN());
   DFF_X1 \buffer_reg[7][4][2][8]  (.D(\input_filter[4][2] [8]), .CK(n_53_7), 
      .Q(\buffer[7][4][2] [8]), .QN());
   DFF_X1 \buffer_reg[7][4][2][7]  (.D(\input_filter[4][2] [7]), .CK(n_53_7), 
      .Q(\buffer[7][4][2] [7]), .QN());
   DFF_X1 \buffer_reg[7][4][2][6]  (.D(\input_filter[4][2] [6]), .CK(n_53_7), 
      .Q(\buffer[7][4][2] [6]), .QN());
   DFF_X1 \buffer_reg[7][4][2][5]  (.D(\input_filter[4][2] [5]), .CK(n_53_7), 
      .Q(\buffer[7][4][2] [5]), .QN());
   DFF_X1 \buffer_reg[7][4][2][4]  (.D(\input_filter[4][2] [4]), .CK(n_53_7), 
      .Q(\buffer[7][4][2] [4]), .QN());
   DFF_X1 \buffer_reg[7][4][2][3]  (.D(\input_filter[4][2] [3]), .CK(n_53_7), 
      .Q(\buffer[7][4][2] [3]), .QN());
   DFF_X1 \buffer_reg[7][4][2][2]  (.D(\input_filter[4][2] [2]), .CK(n_53_7), 
      .Q(\buffer[7][4][2] [2]), .QN());
   DFF_X1 \buffer_reg[7][4][2][1]  (.D(\input_filter[4][2] [1]), .CK(n_53_7), 
      .Q(\buffer[7][4][2] [1]), .QN());
   DFF_X1 \buffer_reg[7][4][2][0]  (.D(\input_filter[4][2] [0]), .CK(n_53_7), 
      .Q(\buffer[7][4][2] [0]), .QN());
   DFF_X1 \buffer_reg[6][4][2][15]  (.D(\input_filter[4][2] [15]), .CK(n_53_6), 
      .Q(\buffer[6][4][2] [15]), .QN());
   DFF_X1 \buffer_reg[6][4][2][14]  (.D(\input_filter[4][2] [14]), .CK(n_53_6), 
      .Q(\buffer[6][4][2] [14]), .QN());
   DFF_X1 \buffer_reg[6][4][2][13]  (.D(\input_filter[4][2] [13]), .CK(n_53_6), 
      .Q(\buffer[6][4][2] [13]), .QN());
   DFF_X1 \buffer_reg[6][4][2][12]  (.D(\input_filter[4][2] [12]), .CK(n_53_6), 
      .Q(\buffer[6][4][2] [12]), .QN());
   DFF_X1 \buffer_reg[6][4][2][11]  (.D(\input_filter[4][2] [11]), .CK(n_53_6), 
      .Q(\buffer[6][4][2] [11]), .QN());
   DFF_X1 \buffer_reg[6][4][2][10]  (.D(\input_filter[4][2] [10]), .CK(n_53_6), 
      .Q(\buffer[6][4][2] [10]), .QN());
   DFF_X1 \buffer_reg[6][4][2][9]  (.D(\input_filter[4][2] [9]), .CK(n_53_6), 
      .Q(\buffer[6][4][2] [9]), .QN());
   DFF_X1 \buffer_reg[6][4][2][8]  (.D(\input_filter[4][2] [8]), .CK(n_53_6), 
      .Q(\buffer[6][4][2] [8]), .QN());
   DFF_X1 \buffer_reg[6][4][2][7]  (.D(\input_filter[4][2] [7]), .CK(n_53_6), 
      .Q(\buffer[6][4][2] [7]), .QN());
   DFF_X1 \buffer_reg[6][4][2][6]  (.D(\input_filter[4][2] [6]), .CK(n_53_6), 
      .Q(\buffer[6][4][2] [6]), .QN());
   DFF_X1 \buffer_reg[6][4][2][5]  (.D(\input_filter[4][2] [5]), .CK(n_53_6), 
      .Q(\buffer[6][4][2] [5]), .QN());
   DFF_X1 \buffer_reg[6][4][2][4]  (.D(\input_filter[4][2] [4]), .CK(n_53_6), 
      .Q(\buffer[6][4][2] [4]), .QN());
   DFF_X1 \buffer_reg[6][4][2][3]  (.D(\input_filter[4][2] [3]), .CK(n_53_6), 
      .Q(\buffer[6][4][2] [3]), .QN());
   DFF_X1 \buffer_reg[6][4][2][2]  (.D(\input_filter[4][2] [2]), .CK(n_53_6), 
      .Q(\buffer[6][4][2] [2]), .QN());
   DFF_X1 \buffer_reg[6][4][2][1]  (.D(\input_filter[4][2] [1]), .CK(n_53_6), 
      .Q(\buffer[6][4][2] [1]), .QN());
   DFF_X1 \buffer_reg[6][4][2][0]  (.D(\input_filter[4][2] [0]), .CK(n_53_6), 
      .Q(\buffer[6][4][2] [0]), .QN());
   DFF_X1 \buffer_reg[5][4][2][15]  (.D(\input_filter[4][2] [15]), .CK(n_53_5), 
      .Q(\buffer[5][4][2] [15]), .QN());
   DFF_X1 \buffer_reg[5][4][2][14]  (.D(\input_filter[4][2] [14]), .CK(n_53_5), 
      .Q(\buffer[5][4][2] [14]), .QN());
   DFF_X1 \buffer_reg[5][4][2][13]  (.D(\input_filter[4][2] [13]), .CK(n_53_5), 
      .Q(\buffer[5][4][2] [13]), .QN());
   DFF_X1 \buffer_reg[5][4][2][12]  (.D(\input_filter[4][2] [12]), .CK(n_53_5), 
      .Q(\buffer[5][4][2] [12]), .QN());
   DFF_X1 \buffer_reg[5][4][2][11]  (.D(\input_filter[4][2] [11]), .CK(n_53_5), 
      .Q(\buffer[5][4][2] [11]), .QN());
   DFF_X1 \buffer_reg[5][4][2][10]  (.D(\input_filter[4][2] [10]), .CK(n_53_5), 
      .Q(\buffer[5][4][2] [10]), .QN());
   DFF_X1 \buffer_reg[5][4][2][9]  (.D(\input_filter[4][2] [9]), .CK(n_53_5), 
      .Q(\buffer[5][4][2] [9]), .QN());
   DFF_X1 \buffer_reg[5][4][2][8]  (.D(\input_filter[4][2] [8]), .CK(n_53_5), 
      .Q(\buffer[5][4][2] [8]), .QN());
   DFF_X1 \buffer_reg[5][4][2][7]  (.D(\input_filter[4][2] [7]), .CK(n_53_5), 
      .Q(\buffer[5][4][2] [7]), .QN());
   DFF_X1 \buffer_reg[5][4][2][6]  (.D(\input_filter[4][2] [6]), .CK(n_53_5), 
      .Q(\buffer[5][4][2] [6]), .QN());
   DFF_X1 \buffer_reg[5][4][2][5]  (.D(\input_filter[4][2] [5]), .CK(n_53_5), 
      .Q(\buffer[5][4][2] [5]), .QN());
   DFF_X1 \buffer_reg[5][4][2][4]  (.D(\input_filter[4][2] [4]), .CK(n_53_5), 
      .Q(\buffer[5][4][2] [4]), .QN());
   DFF_X1 \buffer_reg[5][4][2][3]  (.D(\input_filter[4][2] [3]), .CK(n_53_5), 
      .Q(\buffer[5][4][2] [3]), .QN());
   DFF_X1 \buffer_reg[5][4][2][2]  (.D(\input_filter[4][2] [2]), .CK(n_53_5), 
      .Q(\buffer[5][4][2] [2]), .QN());
   DFF_X1 \buffer_reg[5][4][2][1]  (.D(\input_filter[4][2] [1]), .CK(n_53_5), 
      .Q(\buffer[5][4][2] [1]), .QN());
   DFF_X1 \buffer_reg[5][4][2][0]  (.D(\input_filter[4][2] [0]), .CK(n_53_5), 
      .Q(\buffer[5][4][2] [0]), .QN());
   DFF_X1 \buffer_reg[4][4][2][15]  (.D(\input_filter[4][2] [15]), .CK(n_53_4), 
      .Q(\buffer[4][4][2] [15]), .QN());
   DFF_X1 \buffer_reg[4][4][2][14]  (.D(\input_filter[4][2] [14]), .CK(n_53_4), 
      .Q(\buffer[4][4][2] [14]), .QN());
   DFF_X1 \buffer_reg[4][4][2][13]  (.D(\input_filter[4][2] [13]), .CK(n_53_4), 
      .Q(\buffer[4][4][2] [13]), .QN());
   DFF_X1 \buffer_reg[4][4][2][12]  (.D(\input_filter[4][2] [12]), .CK(n_53_4), 
      .Q(\buffer[4][4][2] [12]), .QN());
   DFF_X1 \buffer_reg[4][4][2][11]  (.D(\input_filter[4][2] [11]), .CK(n_53_4), 
      .Q(\buffer[4][4][2] [11]), .QN());
   DFF_X1 \buffer_reg[4][4][2][10]  (.D(\input_filter[4][2] [10]), .CK(n_53_4), 
      .Q(\buffer[4][4][2] [10]), .QN());
   DFF_X1 \buffer_reg[4][4][2][9]  (.D(\input_filter[4][2] [9]), .CK(n_53_4), 
      .Q(\buffer[4][4][2] [9]), .QN());
   DFF_X1 \buffer_reg[4][4][2][8]  (.D(\input_filter[4][2] [8]), .CK(n_53_4), 
      .Q(\buffer[4][4][2] [8]), .QN());
   DFF_X1 \buffer_reg[4][4][2][7]  (.D(\input_filter[4][2] [7]), .CK(n_53_4), 
      .Q(\buffer[4][4][2] [7]), .QN());
   DFF_X1 \buffer_reg[4][4][2][6]  (.D(\input_filter[4][2] [6]), .CK(n_53_4), 
      .Q(\buffer[4][4][2] [6]), .QN());
   DFF_X1 \buffer_reg[4][4][2][5]  (.D(\input_filter[4][2] [5]), .CK(n_53_4), 
      .Q(\buffer[4][4][2] [5]), .QN());
   DFF_X1 \buffer_reg[4][4][2][4]  (.D(\input_filter[4][2] [4]), .CK(n_53_4), 
      .Q(\buffer[4][4][2] [4]), .QN());
   DFF_X1 \buffer_reg[4][4][2][3]  (.D(\input_filter[4][2] [3]), .CK(n_53_4), 
      .Q(\buffer[4][4][2] [3]), .QN());
   DFF_X1 \buffer_reg[4][4][2][2]  (.D(\input_filter[4][2] [2]), .CK(n_53_4), 
      .Q(\buffer[4][4][2] [2]), .QN());
   DFF_X1 \buffer_reg[4][4][2][1]  (.D(\input_filter[4][2] [1]), .CK(n_53_4), 
      .Q(\buffer[4][4][2] [1]), .QN());
   DFF_X1 \buffer_reg[4][4][2][0]  (.D(\input_filter[4][2] [0]), .CK(n_53_4), 
      .Q(\buffer[4][4][2] [0]), .QN());
   DFF_X1 \buffer_reg[3][4][2][15]  (.D(\input_filter[4][2] [15]), .CK(n_53_3), 
      .Q(\buffer[3][4][2] [15]), .QN());
   DFF_X1 \buffer_reg[3][4][2][14]  (.D(\input_filter[4][2] [14]), .CK(n_53_3), 
      .Q(\buffer[3][4][2] [14]), .QN());
   DFF_X1 \buffer_reg[3][4][2][13]  (.D(\input_filter[4][2] [13]), .CK(n_53_3), 
      .Q(\buffer[3][4][2] [13]), .QN());
   DFF_X1 \buffer_reg[3][4][2][12]  (.D(\input_filter[4][2] [12]), .CK(n_53_3), 
      .Q(\buffer[3][4][2] [12]), .QN());
   DFF_X1 \buffer_reg[3][4][2][11]  (.D(\input_filter[4][2] [11]), .CK(n_53_3), 
      .Q(\buffer[3][4][2] [11]), .QN());
   DFF_X1 \buffer_reg[3][4][2][10]  (.D(\input_filter[4][2] [10]), .CK(n_53_3), 
      .Q(\buffer[3][4][2] [10]), .QN());
   DFF_X1 \buffer_reg[3][4][2][9]  (.D(\input_filter[4][2] [9]), .CK(n_53_3), 
      .Q(\buffer[3][4][2] [9]), .QN());
   DFF_X1 \buffer_reg[3][4][2][8]  (.D(\input_filter[4][2] [8]), .CK(n_53_3), 
      .Q(\buffer[3][4][2] [8]), .QN());
   DFF_X1 \buffer_reg[3][4][2][7]  (.D(\input_filter[4][2] [7]), .CK(n_53_3), 
      .Q(\buffer[3][4][2] [7]), .QN());
   DFF_X1 \buffer_reg[3][4][2][6]  (.D(\input_filter[4][2] [6]), .CK(n_53_3), 
      .Q(\buffer[3][4][2] [6]), .QN());
   DFF_X1 \buffer_reg[3][4][2][5]  (.D(\input_filter[4][2] [5]), .CK(n_53_3), 
      .Q(\buffer[3][4][2] [5]), .QN());
   DFF_X1 \buffer_reg[3][4][2][4]  (.D(\input_filter[4][2] [4]), .CK(n_53_3), 
      .Q(\buffer[3][4][2] [4]), .QN());
   DFF_X1 \buffer_reg[3][4][2][3]  (.D(\input_filter[4][2] [3]), .CK(n_53_3), 
      .Q(\buffer[3][4][2] [3]), .QN());
   DFF_X1 \buffer_reg[3][4][2][2]  (.D(\input_filter[4][2] [2]), .CK(n_53_3), 
      .Q(\buffer[3][4][2] [2]), .QN());
   DFF_X1 \buffer_reg[3][4][2][1]  (.D(\input_filter[4][2] [1]), .CK(n_53_3), 
      .Q(\buffer[3][4][2] [1]), .QN());
   DFF_X1 \buffer_reg[3][4][2][0]  (.D(\input_filter[4][2] [0]), .CK(n_53_3), 
      .Q(\buffer[3][4][2] [0]), .QN());
   DFF_X1 \buffer_reg[2][4][2][15]  (.D(\input_filter[4][2] [15]), .CK(n_53_2), 
      .Q(\buffer[2][4][2] [15]), .QN());
   DFF_X1 \buffer_reg[2][4][2][14]  (.D(\input_filter[4][2] [14]), .CK(n_53_2), 
      .Q(\buffer[2][4][2] [14]), .QN());
   DFF_X1 \buffer_reg[2][4][2][13]  (.D(\input_filter[4][2] [13]), .CK(n_53_2), 
      .Q(\buffer[2][4][2] [13]), .QN());
   DFF_X1 \buffer_reg[2][4][2][12]  (.D(\input_filter[4][2] [12]), .CK(n_53_2), 
      .Q(\buffer[2][4][2] [12]), .QN());
   DFF_X1 \buffer_reg[2][4][2][11]  (.D(\input_filter[4][2] [11]), .CK(n_53_2), 
      .Q(\buffer[2][4][2] [11]), .QN());
   DFF_X1 \buffer_reg[2][4][2][10]  (.D(\input_filter[4][2] [10]), .CK(n_53_2), 
      .Q(\buffer[2][4][2] [10]), .QN());
   DFF_X1 \buffer_reg[2][4][2][9]  (.D(\input_filter[4][2] [9]), .CK(n_53_2), 
      .Q(\buffer[2][4][2] [9]), .QN());
   DFF_X1 \buffer_reg[2][4][2][8]  (.D(\input_filter[4][2] [8]), .CK(n_53_2), 
      .Q(\buffer[2][4][2] [8]), .QN());
   DFF_X1 \buffer_reg[2][4][2][7]  (.D(\input_filter[4][2] [7]), .CK(n_53_2), 
      .Q(\buffer[2][4][2] [7]), .QN());
   DFF_X1 \buffer_reg[2][4][2][6]  (.D(\input_filter[4][2] [6]), .CK(n_53_2), 
      .Q(\buffer[2][4][2] [6]), .QN());
   DFF_X1 \buffer_reg[2][4][2][5]  (.D(\input_filter[4][2] [5]), .CK(n_53_2), 
      .Q(\buffer[2][4][2] [5]), .QN());
   DFF_X1 \buffer_reg[2][4][2][4]  (.D(\input_filter[4][2] [4]), .CK(n_53_2), 
      .Q(\buffer[2][4][2] [4]), .QN());
   DFF_X1 \buffer_reg[2][4][2][3]  (.D(\input_filter[4][2] [3]), .CK(n_53_2), 
      .Q(\buffer[2][4][2] [3]), .QN());
   DFF_X1 \buffer_reg[2][4][2][2]  (.D(\input_filter[4][2] [2]), .CK(n_53_2), 
      .Q(\buffer[2][4][2] [2]), .QN());
   DFF_X1 \buffer_reg[2][4][2][1]  (.D(\input_filter[4][2] [1]), .CK(n_53_2), 
      .Q(\buffer[2][4][2] [1]), .QN());
   DFF_X1 \buffer_reg[2][4][2][0]  (.D(\input_filter[4][2] [0]), .CK(n_53_2), 
      .Q(\buffer[2][4][2] [0]), .QN());
   DFF_X1 \buffer_reg[1][4][2][15]  (.D(\input_filter[4][2] [15]), .CK(n_53_1), 
      .Q(\buffer[1][4][2] [15]), .QN());
   DFF_X1 \buffer_reg[1][4][2][14]  (.D(\input_filter[4][2] [14]), .CK(n_53_1), 
      .Q(\buffer[1][4][2] [14]), .QN());
   DFF_X1 \buffer_reg[1][4][2][13]  (.D(\input_filter[4][2] [13]), .CK(n_53_1), 
      .Q(\buffer[1][4][2] [13]), .QN());
   DFF_X1 \buffer_reg[1][4][2][12]  (.D(\input_filter[4][2] [12]), .CK(n_53_1), 
      .Q(\buffer[1][4][2] [12]), .QN());
   DFF_X1 \buffer_reg[1][4][2][11]  (.D(\input_filter[4][2] [11]), .CK(n_53_1), 
      .Q(\buffer[1][4][2] [11]), .QN());
   DFF_X1 \buffer_reg[1][4][2][10]  (.D(\input_filter[4][2] [10]), .CK(n_53_1), 
      .Q(\buffer[1][4][2] [10]), .QN());
   DFF_X1 \buffer_reg[1][4][2][9]  (.D(\input_filter[4][2] [9]), .CK(n_53_1), 
      .Q(\buffer[1][4][2] [9]), .QN());
   DFF_X1 \buffer_reg[1][4][2][8]  (.D(\input_filter[4][2] [8]), .CK(n_53_1), 
      .Q(\buffer[1][4][2] [8]), .QN());
   DFF_X1 \buffer_reg[1][4][2][7]  (.D(\input_filter[4][2] [7]), .CK(n_53_1), 
      .Q(\buffer[1][4][2] [7]), .QN());
   DFF_X1 \buffer_reg[1][4][2][6]  (.D(\input_filter[4][2] [6]), .CK(n_53_1), 
      .Q(\buffer[1][4][2] [6]), .QN());
   DFF_X1 \buffer_reg[1][4][2][5]  (.D(\input_filter[4][2] [5]), .CK(n_53_1), 
      .Q(\buffer[1][4][2] [5]), .QN());
   DFF_X1 \buffer_reg[1][4][2][4]  (.D(\input_filter[4][2] [4]), .CK(n_53_1), 
      .Q(\buffer[1][4][2] [4]), .QN());
   DFF_X1 \buffer_reg[1][4][2][3]  (.D(\input_filter[4][2] [3]), .CK(n_53_1), 
      .Q(\buffer[1][4][2] [3]), .QN());
   DFF_X1 \buffer_reg[1][4][2][2]  (.D(\input_filter[4][2] [2]), .CK(n_53_1), 
      .Q(\buffer[1][4][2] [2]), .QN());
   DFF_X1 \buffer_reg[1][4][2][1]  (.D(\input_filter[4][2] [1]), .CK(n_53_1), 
      .Q(\buffer[1][4][2] [1]), .QN());
   DFF_X1 \buffer_reg[1][4][2][0]  (.D(\input_filter[4][2] [0]), .CK(n_53_1), 
      .Q(\buffer[1][4][2] [0]), .QN());
   DFF_X1 \buffer_reg[0][4][2][15]  (.D(\input_filter[4][2] [15]), .CK(n_53_0), 
      .Q(\buffer[0][4][2] [15]), .QN());
   DFF_X1 \buffer_reg[0][4][2][14]  (.D(\input_filter[4][2] [14]), .CK(n_53_0), 
      .Q(\buffer[0][4][2] [14]), .QN());
   DFF_X1 \buffer_reg[0][4][2][13]  (.D(\input_filter[4][2] [13]), .CK(n_53_0), 
      .Q(\buffer[0][4][2] [13]), .QN());
   DFF_X1 \buffer_reg[0][4][2][12]  (.D(\input_filter[4][2] [12]), .CK(n_53_0), 
      .Q(\buffer[0][4][2] [12]), .QN());
   DFF_X1 \buffer_reg[0][4][2][11]  (.D(\input_filter[4][2] [11]), .CK(n_53_0), 
      .Q(\buffer[0][4][2] [11]), .QN());
   DFF_X1 \buffer_reg[0][4][2][10]  (.D(\input_filter[4][2] [10]), .CK(n_53_0), 
      .Q(\buffer[0][4][2] [10]), .QN());
   DFF_X1 \buffer_reg[0][4][2][9]  (.D(\input_filter[4][2] [9]), .CK(n_53_0), 
      .Q(\buffer[0][4][2] [9]), .QN());
   DFF_X1 \buffer_reg[0][4][2][8]  (.D(\input_filter[4][2] [8]), .CK(n_53_0), 
      .Q(\buffer[0][4][2] [8]), .QN());
   DFF_X1 \buffer_reg[0][4][2][7]  (.D(\input_filter[4][2] [7]), .CK(n_53_0), 
      .Q(\buffer[0][4][2] [7]), .QN());
   DFF_X1 \buffer_reg[0][4][2][6]  (.D(\input_filter[4][2] [6]), .CK(n_53_0), 
      .Q(\buffer[0][4][2] [6]), .QN());
   DFF_X1 \buffer_reg[0][4][2][5]  (.D(\input_filter[4][2] [5]), .CK(n_53_0), 
      .Q(\buffer[0][4][2] [5]), .QN());
   DFF_X1 \buffer_reg[0][4][2][4]  (.D(\input_filter[4][2] [4]), .CK(n_53_0), 
      .Q(\buffer[0][4][2] [4]), .QN());
   DFF_X1 \buffer_reg[0][4][2][3]  (.D(\input_filter[4][2] [3]), .CK(n_53_0), 
      .Q(\buffer[0][4][2] [3]), .QN());
   DFF_X1 \buffer_reg[0][4][2][2]  (.D(\input_filter[4][2] [2]), .CK(n_53_0), 
      .Q(\buffer[0][4][2] [2]), .QN());
   DFF_X1 \buffer_reg[0][4][2][1]  (.D(\input_filter[4][2] [1]), .CK(n_53_0), 
      .Q(\buffer[0][4][2] [1]), .QN());
   DFF_X1 \buffer_reg[0][4][2][0]  (.D(\input_filter[4][2] [0]), .CK(n_53_0), 
      .Q(\buffer[0][4][2] [0]), .QN());
   DFF_X1 \buffer_reg[15][4][1][15]  (.D(\input_filter[4][1] [15]), .CK(n_53_15), 
      .Q(\buffer[15][4][1] [15]), .QN());
   DFF_X1 \buffer_reg[15][4][1][14]  (.D(\input_filter[4][1] [14]), .CK(n_53_15), 
      .Q(\buffer[15][4][1] [14]), .QN());
   DFF_X1 \buffer_reg[15][4][1][13]  (.D(\input_filter[4][1] [13]), .CK(n_53_15), 
      .Q(\buffer[15][4][1] [13]), .QN());
   DFF_X1 \buffer_reg[15][4][1][12]  (.D(\input_filter[4][1] [12]), .CK(n_53_15), 
      .Q(\buffer[15][4][1] [12]), .QN());
   DFF_X1 \buffer_reg[15][4][1][11]  (.D(\input_filter[4][1] [11]), .CK(n_53_15), 
      .Q(\buffer[15][4][1] [11]), .QN());
   DFF_X1 \buffer_reg[15][4][1][10]  (.D(\input_filter[4][1] [10]), .CK(n_53_15), 
      .Q(\buffer[15][4][1] [10]), .QN());
   DFF_X1 \buffer_reg[15][4][1][9]  (.D(\input_filter[4][1] [9]), .CK(n_53_15), 
      .Q(\buffer[15][4][1] [9]), .QN());
   DFF_X1 \buffer_reg[15][4][1][8]  (.D(\input_filter[4][1] [8]), .CK(n_53_15), 
      .Q(\buffer[15][4][1] [8]), .QN());
   DFF_X1 \buffer_reg[15][4][1][7]  (.D(\input_filter[4][1] [7]), .CK(n_53_15), 
      .Q(\buffer[15][4][1] [7]), .QN());
   DFF_X1 \buffer_reg[15][4][1][6]  (.D(\input_filter[4][1] [6]), .CK(n_53_15), 
      .Q(\buffer[15][4][1] [6]), .QN());
   DFF_X1 \buffer_reg[15][4][1][5]  (.D(\input_filter[4][1] [5]), .CK(n_53_15), 
      .Q(\buffer[15][4][1] [5]), .QN());
   DFF_X1 \buffer_reg[15][4][1][4]  (.D(\input_filter[4][1] [4]), .CK(n_53_15), 
      .Q(\buffer[15][4][1] [4]), .QN());
   DFF_X1 \buffer_reg[15][4][1][3]  (.D(\input_filter[4][1] [3]), .CK(n_53_15), 
      .Q(\buffer[15][4][1] [3]), .QN());
   DFF_X1 \buffer_reg[15][4][1][2]  (.D(\input_filter[4][1] [2]), .CK(n_53_15), 
      .Q(\buffer[15][4][1] [2]), .QN());
   DFF_X1 \buffer_reg[15][4][1][1]  (.D(\input_filter[4][1] [1]), .CK(n_53_15), 
      .Q(\buffer[15][4][1] [1]), .QN());
   DFF_X1 \buffer_reg[15][4][1][0]  (.D(\input_filter[4][1] [0]), .CK(n_53_15), 
      .Q(\buffer[15][4][1] [0]), .QN());
   DFF_X1 \buffer_reg[14][4][1][15]  (.D(\input_filter[4][1] [15]), .CK(n_53_14), 
      .Q(\buffer[14][4][1] [15]), .QN());
   DFF_X1 \buffer_reg[14][4][1][14]  (.D(\input_filter[4][1] [14]), .CK(n_53_14), 
      .Q(\buffer[14][4][1] [14]), .QN());
   DFF_X1 \buffer_reg[14][4][1][13]  (.D(\input_filter[4][1] [13]), .CK(n_53_14), 
      .Q(\buffer[14][4][1] [13]), .QN());
   DFF_X1 \buffer_reg[14][4][1][12]  (.D(\input_filter[4][1] [12]), .CK(n_53_14), 
      .Q(\buffer[14][4][1] [12]), .QN());
   DFF_X1 \buffer_reg[14][4][1][11]  (.D(\input_filter[4][1] [11]), .CK(n_53_14), 
      .Q(\buffer[14][4][1] [11]), .QN());
   DFF_X1 \buffer_reg[14][4][1][10]  (.D(\input_filter[4][1] [10]), .CK(n_53_14), 
      .Q(\buffer[14][4][1] [10]), .QN());
   DFF_X1 \buffer_reg[14][4][1][9]  (.D(\input_filter[4][1] [9]), .CK(n_53_14), 
      .Q(\buffer[14][4][1] [9]), .QN());
   DFF_X1 \buffer_reg[14][4][1][8]  (.D(\input_filter[4][1] [8]), .CK(n_53_14), 
      .Q(\buffer[14][4][1] [8]), .QN());
   DFF_X1 \buffer_reg[14][4][1][7]  (.D(\input_filter[4][1] [7]), .CK(n_53_14), 
      .Q(\buffer[14][4][1] [7]), .QN());
   DFF_X1 \buffer_reg[14][4][1][6]  (.D(\input_filter[4][1] [6]), .CK(n_53_14), 
      .Q(\buffer[14][4][1] [6]), .QN());
   DFF_X1 \buffer_reg[14][4][1][5]  (.D(\input_filter[4][1] [5]), .CK(n_53_14), 
      .Q(\buffer[14][4][1] [5]), .QN());
   DFF_X1 \buffer_reg[14][4][1][4]  (.D(\input_filter[4][1] [4]), .CK(n_53_14), 
      .Q(\buffer[14][4][1] [4]), .QN());
   DFF_X1 \buffer_reg[14][4][1][3]  (.D(\input_filter[4][1] [3]), .CK(n_53_14), 
      .Q(\buffer[14][4][1] [3]), .QN());
   DFF_X1 \buffer_reg[14][4][1][2]  (.D(\input_filter[4][1] [2]), .CK(n_53_14), 
      .Q(\buffer[14][4][1] [2]), .QN());
   DFF_X1 \buffer_reg[14][4][1][1]  (.D(\input_filter[4][1] [1]), .CK(n_53_14), 
      .Q(\buffer[14][4][1] [1]), .QN());
   DFF_X1 \buffer_reg[14][4][1][0]  (.D(\input_filter[4][1] [0]), .CK(n_53_14), 
      .Q(\buffer[14][4][1] [0]), .QN());
   DFF_X1 \buffer_reg[13][4][1][15]  (.D(\input_filter[4][1] [15]), .CK(n_53_13), 
      .Q(\buffer[13][4][1] [15]), .QN());
   DFF_X1 \buffer_reg[13][4][1][14]  (.D(\input_filter[4][1] [14]), .CK(n_53_13), 
      .Q(\buffer[13][4][1] [14]), .QN());
   DFF_X1 \buffer_reg[13][4][1][13]  (.D(\input_filter[4][1] [13]), .CK(n_53_13), 
      .Q(\buffer[13][4][1] [13]), .QN());
   DFF_X1 \buffer_reg[13][4][1][12]  (.D(\input_filter[4][1] [12]), .CK(n_53_13), 
      .Q(\buffer[13][4][1] [12]), .QN());
   DFF_X1 \buffer_reg[13][4][1][11]  (.D(\input_filter[4][1] [11]), .CK(n_53_13), 
      .Q(\buffer[13][4][1] [11]), .QN());
   DFF_X1 \buffer_reg[13][4][1][10]  (.D(\input_filter[4][1] [10]), .CK(n_53_13), 
      .Q(\buffer[13][4][1] [10]), .QN());
   DFF_X1 \buffer_reg[13][4][1][9]  (.D(\input_filter[4][1] [9]), .CK(n_53_13), 
      .Q(\buffer[13][4][1] [9]), .QN());
   DFF_X1 \buffer_reg[13][4][1][8]  (.D(\input_filter[4][1] [8]), .CK(n_53_13), 
      .Q(\buffer[13][4][1] [8]), .QN());
   DFF_X1 \buffer_reg[13][4][1][7]  (.D(\input_filter[4][1] [7]), .CK(n_53_13), 
      .Q(\buffer[13][4][1] [7]), .QN());
   DFF_X1 \buffer_reg[13][4][1][6]  (.D(\input_filter[4][1] [6]), .CK(n_53_13), 
      .Q(\buffer[13][4][1] [6]), .QN());
   DFF_X1 \buffer_reg[13][4][1][5]  (.D(\input_filter[4][1] [5]), .CK(n_53_13), 
      .Q(\buffer[13][4][1] [5]), .QN());
   DFF_X1 \buffer_reg[13][4][1][4]  (.D(\input_filter[4][1] [4]), .CK(n_53_13), 
      .Q(\buffer[13][4][1] [4]), .QN());
   DFF_X1 \buffer_reg[13][4][1][3]  (.D(\input_filter[4][1] [3]), .CK(n_53_13), 
      .Q(\buffer[13][4][1] [3]), .QN());
   DFF_X1 \buffer_reg[13][4][1][2]  (.D(\input_filter[4][1] [2]), .CK(n_53_13), 
      .Q(\buffer[13][4][1] [2]), .QN());
   DFF_X1 \buffer_reg[13][4][1][1]  (.D(\input_filter[4][1] [1]), .CK(n_53_13), 
      .Q(\buffer[13][4][1] [1]), .QN());
   DFF_X1 \buffer_reg[13][4][1][0]  (.D(\input_filter[4][1] [0]), .CK(n_53_13), 
      .Q(\buffer[13][4][1] [0]), .QN());
   DFF_X1 \buffer_reg[12][4][1][15]  (.D(\input_filter[4][1] [15]), .CK(n_53_12), 
      .Q(\buffer[12][4][1] [15]), .QN());
   DFF_X1 \buffer_reg[12][4][1][14]  (.D(\input_filter[4][1] [14]), .CK(n_53_12), 
      .Q(\buffer[12][4][1] [14]), .QN());
   DFF_X1 \buffer_reg[12][4][1][13]  (.D(\input_filter[4][1] [13]), .CK(n_53_12), 
      .Q(\buffer[12][4][1] [13]), .QN());
   DFF_X1 \buffer_reg[12][4][1][12]  (.D(\input_filter[4][1] [12]), .CK(n_53_12), 
      .Q(\buffer[12][4][1] [12]), .QN());
   DFF_X1 \buffer_reg[12][4][1][11]  (.D(\input_filter[4][1] [11]), .CK(n_53_12), 
      .Q(\buffer[12][4][1] [11]), .QN());
   DFF_X1 \buffer_reg[12][4][1][10]  (.D(\input_filter[4][1] [10]), .CK(n_53_12), 
      .Q(\buffer[12][4][1] [10]), .QN());
   DFF_X1 \buffer_reg[12][4][1][9]  (.D(\input_filter[4][1] [9]), .CK(n_53_12), 
      .Q(\buffer[12][4][1] [9]), .QN());
   DFF_X1 \buffer_reg[12][4][1][8]  (.D(\input_filter[4][1] [8]), .CK(n_53_12), 
      .Q(\buffer[12][4][1] [8]), .QN());
   DFF_X1 \buffer_reg[12][4][1][7]  (.D(\input_filter[4][1] [7]), .CK(n_53_12), 
      .Q(\buffer[12][4][1] [7]), .QN());
   DFF_X1 \buffer_reg[12][4][1][6]  (.D(\input_filter[4][1] [6]), .CK(n_53_12), 
      .Q(\buffer[12][4][1] [6]), .QN());
   DFF_X1 \buffer_reg[12][4][1][5]  (.D(\input_filter[4][1] [5]), .CK(n_53_12), 
      .Q(\buffer[12][4][1] [5]), .QN());
   DFF_X1 \buffer_reg[12][4][1][4]  (.D(\input_filter[4][1] [4]), .CK(n_53_12), 
      .Q(\buffer[12][4][1] [4]), .QN());
   DFF_X1 \buffer_reg[12][4][1][3]  (.D(\input_filter[4][1] [3]), .CK(n_53_12), 
      .Q(\buffer[12][4][1] [3]), .QN());
   DFF_X1 \buffer_reg[12][4][1][2]  (.D(\input_filter[4][1] [2]), .CK(n_53_12), 
      .Q(\buffer[12][4][1] [2]), .QN());
   DFF_X1 \buffer_reg[12][4][1][1]  (.D(\input_filter[4][1] [1]), .CK(n_53_12), 
      .Q(\buffer[12][4][1] [1]), .QN());
   DFF_X1 \buffer_reg[12][4][1][0]  (.D(\input_filter[4][1] [0]), .CK(n_53_12), 
      .Q(\buffer[12][4][1] [0]), .QN());
   DFF_X1 \buffer_reg[11][4][1][15]  (.D(\input_filter[4][1] [15]), .CK(n_53_11), 
      .Q(\buffer[11][4][1] [15]), .QN());
   DFF_X1 \buffer_reg[11][4][1][14]  (.D(\input_filter[4][1] [14]), .CK(n_53_11), 
      .Q(\buffer[11][4][1] [14]), .QN());
   DFF_X1 \buffer_reg[11][4][1][13]  (.D(\input_filter[4][1] [13]), .CK(n_53_11), 
      .Q(\buffer[11][4][1] [13]), .QN());
   DFF_X1 \buffer_reg[11][4][1][12]  (.D(\input_filter[4][1] [12]), .CK(n_53_11), 
      .Q(\buffer[11][4][1] [12]), .QN());
   DFF_X1 \buffer_reg[11][4][1][11]  (.D(\input_filter[4][1] [11]), .CK(n_53_11), 
      .Q(\buffer[11][4][1] [11]), .QN());
   DFF_X1 \buffer_reg[11][4][1][10]  (.D(\input_filter[4][1] [10]), .CK(n_53_11), 
      .Q(\buffer[11][4][1] [10]), .QN());
   DFF_X1 \buffer_reg[11][4][1][9]  (.D(\input_filter[4][1] [9]), .CK(n_53_11), 
      .Q(\buffer[11][4][1] [9]), .QN());
   DFF_X1 \buffer_reg[11][4][1][8]  (.D(\input_filter[4][1] [8]), .CK(n_53_11), 
      .Q(\buffer[11][4][1] [8]), .QN());
   DFF_X1 \buffer_reg[11][4][1][7]  (.D(\input_filter[4][1] [7]), .CK(n_53_11), 
      .Q(\buffer[11][4][1] [7]), .QN());
   DFF_X1 \buffer_reg[11][4][1][6]  (.D(\input_filter[4][1] [6]), .CK(n_53_11), 
      .Q(\buffer[11][4][1] [6]), .QN());
   DFF_X1 \buffer_reg[11][4][1][5]  (.D(\input_filter[4][1] [5]), .CK(n_53_11), 
      .Q(\buffer[11][4][1] [5]), .QN());
   DFF_X1 \buffer_reg[11][4][1][4]  (.D(\input_filter[4][1] [4]), .CK(n_53_11), 
      .Q(\buffer[11][4][1] [4]), .QN());
   DFF_X1 \buffer_reg[11][4][1][3]  (.D(\input_filter[4][1] [3]), .CK(n_53_11), 
      .Q(\buffer[11][4][1] [3]), .QN());
   DFF_X1 \buffer_reg[11][4][1][2]  (.D(\input_filter[4][1] [2]), .CK(n_53_11), 
      .Q(\buffer[11][4][1] [2]), .QN());
   DFF_X1 \buffer_reg[11][4][1][1]  (.D(\input_filter[4][1] [1]), .CK(n_53_11), 
      .Q(\buffer[11][4][1] [1]), .QN());
   DFF_X1 \buffer_reg[11][4][1][0]  (.D(\input_filter[4][1] [0]), .CK(n_53_11), 
      .Q(\buffer[11][4][1] [0]), .QN());
   DFF_X1 \buffer_reg[10][4][1][15]  (.D(\input_filter[4][1] [15]), .CK(n_53_10), 
      .Q(\buffer[10][4][1] [15]), .QN());
   DFF_X1 \buffer_reg[10][4][1][14]  (.D(\input_filter[4][1] [14]), .CK(n_53_10), 
      .Q(\buffer[10][4][1] [14]), .QN());
   DFF_X1 \buffer_reg[10][4][1][13]  (.D(\input_filter[4][1] [13]), .CK(n_53_10), 
      .Q(\buffer[10][4][1] [13]), .QN());
   DFF_X1 \buffer_reg[10][4][1][12]  (.D(\input_filter[4][1] [12]), .CK(n_53_10), 
      .Q(\buffer[10][4][1] [12]), .QN());
   DFF_X1 \buffer_reg[10][4][1][11]  (.D(\input_filter[4][1] [11]), .CK(n_53_10), 
      .Q(\buffer[10][4][1] [11]), .QN());
   DFF_X1 \buffer_reg[10][4][1][10]  (.D(\input_filter[4][1] [10]), .CK(n_53_10), 
      .Q(\buffer[10][4][1] [10]), .QN());
   DFF_X1 \buffer_reg[10][4][1][9]  (.D(\input_filter[4][1] [9]), .CK(n_53_10), 
      .Q(\buffer[10][4][1] [9]), .QN());
   DFF_X1 \buffer_reg[10][4][1][8]  (.D(\input_filter[4][1] [8]), .CK(n_53_10), 
      .Q(\buffer[10][4][1] [8]), .QN());
   DFF_X1 \buffer_reg[10][4][1][7]  (.D(\input_filter[4][1] [7]), .CK(n_53_10), 
      .Q(\buffer[10][4][1] [7]), .QN());
   DFF_X1 \buffer_reg[10][4][1][6]  (.D(\input_filter[4][1] [6]), .CK(n_53_10), 
      .Q(\buffer[10][4][1] [6]), .QN());
   DFF_X1 \buffer_reg[10][4][1][5]  (.D(\input_filter[4][1] [5]), .CK(n_53_10), 
      .Q(\buffer[10][4][1] [5]), .QN());
   DFF_X1 \buffer_reg[10][4][1][4]  (.D(\input_filter[4][1] [4]), .CK(n_53_10), 
      .Q(\buffer[10][4][1] [4]), .QN());
   DFF_X1 \buffer_reg[10][4][1][3]  (.D(\input_filter[4][1] [3]), .CK(n_53_10), 
      .Q(\buffer[10][4][1] [3]), .QN());
   DFF_X1 \buffer_reg[10][4][1][2]  (.D(\input_filter[4][1] [2]), .CK(n_53_10), 
      .Q(\buffer[10][4][1] [2]), .QN());
   DFF_X1 \buffer_reg[10][4][1][1]  (.D(\input_filter[4][1] [1]), .CK(n_53_10), 
      .Q(\buffer[10][4][1] [1]), .QN());
   DFF_X1 \buffer_reg[10][4][1][0]  (.D(\input_filter[4][1] [0]), .CK(n_53_10), 
      .Q(\buffer[10][4][1] [0]), .QN());
   DFF_X1 \buffer_reg[9][4][1][15]  (.D(\input_filter[4][1] [15]), .CK(n_53_9), 
      .Q(\buffer[9][4][1] [15]), .QN());
   DFF_X1 \buffer_reg[9][4][1][14]  (.D(\input_filter[4][1] [14]), .CK(n_53_9), 
      .Q(\buffer[9][4][1] [14]), .QN());
   DFF_X1 \buffer_reg[9][4][1][13]  (.D(\input_filter[4][1] [13]), .CK(n_53_9), 
      .Q(\buffer[9][4][1] [13]), .QN());
   DFF_X1 \buffer_reg[9][4][1][12]  (.D(\input_filter[4][1] [12]), .CK(n_53_9), 
      .Q(\buffer[9][4][1] [12]), .QN());
   DFF_X1 \buffer_reg[9][4][1][11]  (.D(\input_filter[4][1] [11]), .CK(n_53_9), 
      .Q(\buffer[9][4][1] [11]), .QN());
   DFF_X1 \buffer_reg[9][4][1][10]  (.D(\input_filter[4][1] [10]), .CK(n_53_9), 
      .Q(\buffer[9][4][1] [10]), .QN());
   DFF_X1 \buffer_reg[9][4][1][9]  (.D(\input_filter[4][1] [9]), .CK(n_53_9), 
      .Q(\buffer[9][4][1] [9]), .QN());
   DFF_X1 \buffer_reg[9][4][1][8]  (.D(\input_filter[4][1] [8]), .CK(n_53_9), 
      .Q(\buffer[9][4][1] [8]), .QN());
   DFF_X1 \buffer_reg[9][4][1][7]  (.D(\input_filter[4][1] [7]), .CK(n_53_9), 
      .Q(\buffer[9][4][1] [7]), .QN());
   DFF_X1 \buffer_reg[9][4][1][6]  (.D(\input_filter[4][1] [6]), .CK(n_53_9), 
      .Q(\buffer[9][4][1] [6]), .QN());
   DFF_X1 \buffer_reg[9][4][1][5]  (.D(\input_filter[4][1] [5]), .CK(n_53_9), 
      .Q(\buffer[9][4][1] [5]), .QN());
   DFF_X1 \buffer_reg[9][4][1][4]  (.D(\input_filter[4][1] [4]), .CK(n_53_9), 
      .Q(\buffer[9][4][1] [4]), .QN());
   DFF_X1 \buffer_reg[9][4][1][3]  (.D(\input_filter[4][1] [3]), .CK(n_53_9), 
      .Q(\buffer[9][4][1] [3]), .QN());
   DFF_X1 \buffer_reg[9][4][1][2]  (.D(\input_filter[4][1] [2]), .CK(n_53_9), 
      .Q(\buffer[9][4][1] [2]), .QN());
   DFF_X1 \buffer_reg[9][4][1][1]  (.D(\input_filter[4][1] [1]), .CK(n_53_9), 
      .Q(\buffer[9][4][1] [1]), .QN());
   DFF_X1 \buffer_reg[9][4][1][0]  (.D(\input_filter[4][1] [0]), .CK(n_53_9), 
      .Q(\buffer[9][4][1] [0]), .QN());
   DFF_X1 \buffer_reg[8][4][1][15]  (.D(\input_filter[4][1] [15]), .CK(n_53_8), 
      .Q(\buffer[8][4][1] [15]), .QN());
   DFF_X1 \buffer_reg[8][4][1][14]  (.D(\input_filter[4][1] [14]), .CK(n_53_8), 
      .Q(\buffer[8][4][1] [14]), .QN());
   DFF_X1 \buffer_reg[8][4][1][13]  (.D(\input_filter[4][1] [13]), .CK(n_53_8), 
      .Q(\buffer[8][4][1] [13]), .QN());
   DFF_X1 \buffer_reg[8][4][1][12]  (.D(\input_filter[4][1] [12]), .CK(n_53_8), 
      .Q(\buffer[8][4][1] [12]), .QN());
   DFF_X1 \buffer_reg[8][4][1][11]  (.D(\input_filter[4][1] [11]), .CK(n_53_8), 
      .Q(\buffer[8][4][1] [11]), .QN());
   DFF_X1 \buffer_reg[8][4][1][10]  (.D(\input_filter[4][1] [10]), .CK(n_53_8), 
      .Q(\buffer[8][4][1] [10]), .QN());
   DFF_X1 \buffer_reg[8][4][1][9]  (.D(\input_filter[4][1] [9]), .CK(n_53_8), 
      .Q(\buffer[8][4][1] [9]), .QN());
   DFF_X1 \buffer_reg[8][4][1][8]  (.D(\input_filter[4][1] [8]), .CK(n_53_8), 
      .Q(\buffer[8][4][1] [8]), .QN());
   DFF_X1 \buffer_reg[8][4][1][7]  (.D(\input_filter[4][1] [7]), .CK(n_53_8), 
      .Q(\buffer[8][4][1] [7]), .QN());
   DFF_X1 \buffer_reg[8][4][1][6]  (.D(\input_filter[4][1] [6]), .CK(n_53_8), 
      .Q(\buffer[8][4][1] [6]), .QN());
   DFF_X1 \buffer_reg[8][4][1][5]  (.D(\input_filter[4][1] [5]), .CK(n_53_8), 
      .Q(\buffer[8][4][1] [5]), .QN());
   DFF_X1 \buffer_reg[8][4][1][4]  (.D(\input_filter[4][1] [4]), .CK(n_53_8), 
      .Q(\buffer[8][4][1] [4]), .QN());
   DFF_X1 \buffer_reg[8][4][1][3]  (.D(\input_filter[4][1] [3]), .CK(n_53_8), 
      .Q(\buffer[8][4][1] [3]), .QN());
   DFF_X1 \buffer_reg[8][4][1][2]  (.D(\input_filter[4][1] [2]), .CK(n_53_8), 
      .Q(\buffer[8][4][1] [2]), .QN());
   DFF_X1 \buffer_reg[8][4][1][1]  (.D(\input_filter[4][1] [1]), .CK(n_53_8), 
      .Q(\buffer[8][4][1] [1]), .QN());
   DFF_X1 \buffer_reg[8][4][1][0]  (.D(\input_filter[4][1] [0]), .CK(n_53_8), 
      .Q(\buffer[8][4][1] [0]), .QN());
   DFF_X1 \buffer_reg[7][4][1][15]  (.D(\input_filter[4][1] [15]), .CK(n_53_7), 
      .Q(\buffer[7][4][1] [15]), .QN());
   DFF_X1 \buffer_reg[7][4][1][14]  (.D(\input_filter[4][1] [14]), .CK(n_53_7), 
      .Q(\buffer[7][4][1] [14]), .QN());
   DFF_X1 \buffer_reg[7][4][1][13]  (.D(\input_filter[4][1] [13]), .CK(n_53_7), 
      .Q(\buffer[7][4][1] [13]), .QN());
   DFF_X1 \buffer_reg[7][4][1][12]  (.D(\input_filter[4][1] [12]), .CK(n_53_7), 
      .Q(\buffer[7][4][1] [12]), .QN());
   DFF_X1 \buffer_reg[7][4][1][11]  (.D(\input_filter[4][1] [11]), .CK(n_53_7), 
      .Q(\buffer[7][4][1] [11]), .QN());
   DFF_X1 \buffer_reg[7][4][1][10]  (.D(\input_filter[4][1] [10]), .CK(n_53_7), 
      .Q(\buffer[7][4][1] [10]), .QN());
   DFF_X1 \buffer_reg[7][4][1][9]  (.D(\input_filter[4][1] [9]), .CK(n_53_7), 
      .Q(\buffer[7][4][1] [9]), .QN());
   DFF_X1 \buffer_reg[7][4][1][8]  (.D(\input_filter[4][1] [8]), .CK(n_53_7), 
      .Q(\buffer[7][4][1] [8]), .QN());
   DFF_X1 \buffer_reg[7][4][1][7]  (.D(\input_filter[4][1] [7]), .CK(n_53_7), 
      .Q(\buffer[7][4][1] [7]), .QN());
   DFF_X1 \buffer_reg[7][4][1][6]  (.D(\input_filter[4][1] [6]), .CK(n_53_7), 
      .Q(\buffer[7][4][1] [6]), .QN());
   DFF_X1 \buffer_reg[7][4][1][5]  (.D(\input_filter[4][1] [5]), .CK(n_53_7), 
      .Q(\buffer[7][4][1] [5]), .QN());
   DFF_X1 \buffer_reg[7][4][1][4]  (.D(\input_filter[4][1] [4]), .CK(n_53_7), 
      .Q(\buffer[7][4][1] [4]), .QN());
   DFF_X1 \buffer_reg[7][4][1][3]  (.D(\input_filter[4][1] [3]), .CK(n_53_7), 
      .Q(\buffer[7][4][1] [3]), .QN());
   DFF_X1 \buffer_reg[7][4][1][2]  (.D(\input_filter[4][1] [2]), .CK(n_53_7), 
      .Q(\buffer[7][4][1] [2]), .QN());
   DFF_X1 \buffer_reg[7][4][1][1]  (.D(\input_filter[4][1] [1]), .CK(n_53_7), 
      .Q(\buffer[7][4][1] [1]), .QN());
   DFF_X1 \buffer_reg[7][4][1][0]  (.D(\input_filter[4][1] [0]), .CK(n_53_7), 
      .Q(\buffer[7][4][1] [0]), .QN());
   DFF_X1 \buffer_reg[6][4][1][15]  (.D(\input_filter[4][1] [15]), .CK(n_53_6), 
      .Q(\buffer[6][4][1] [15]), .QN());
   DFF_X1 \buffer_reg[6][4][1][14]  (.D(\input_filter[4][1] [14]), .CK(n_53_6), 
      .Q(\buffer[6][4][1] [14]), .QN());
   DFF_X1 \buffer_reg[6][4][1][13]  (.D(\input_filter[4][1] [13]), .CK(n_53_6), 
      .Q(\buffer[6][4][1] [13]), .QN());
   DFF_X1 \buffer_reg[6][4][1][12]  (.D(\input_filter[4][1] [12]), .CK(n_53_6), 
      .Q(\buffer[6][4][1] [12]), .QN());
   DFF_X1 \buffer_reg[6][4][1][11]  (.D(\input_filter[4][1] [11]), .CK(n_53_6), 
      .Q(\buffer[6][4][1] [11]), .QN());
   DFF_X1 \buffer_reg[6][4][1][10]  (.D(\input_filter[4][1] [10]), .CK(n_53_6), 
      .Q(\buffer[6][4][1] [10]), .QN());
   DFF_X1 \buffer_reg[6][4][1][9]  (.D(\input_filter[4][1] [9]), .CK(n_53_6), 
      .Q(\buffer[6][4][1] [9]), .QN());
   DFF_X1 \buffer_reg[6][4][1][8]  (.D(\input_filter[4][1] [8]), .CK(n_53_6), 
      .Q(\buffer[6][4][1] [8]), .QN());
   DFF_X1 \buffer_reg[6][4][1][7]  (.D(\input_filter[4][1] [7]), .CK(n_53_6), 
      .Q(\buffer[6][4][1] [7]), .QN());
   DFF_X1 \buffer_reg[6][4][1][6]  (.D(\input_filter[4][1] [6]), .CK(n_53_6), 
      .Q(\buffer[6][4][1] [6]), .QN());
   DFF_X1 \buffer_reg[6][4][1][5]  (.D(\input_filter[4][1] [5]), .CK(n_53_6), 
      .Q(\buffer[6][4][1] [5]), .QN());
   DFF_X1 \buffer_reg[6][4][1][4]  (.D(\input_filter[4][1] [4]), .CK(n_53_6), 
      .Q(\buffer[6][4][1] [4]), .QN());
   DFF_X1 \buffer_reg[6][4][1][3]  (.D(\input_filter[4][1] [3]), .CK(n_53_6), 
      .Q(\buffer[6][4][1] [3]), .QN());
   DFF_X1 \buffer_reg[6][4][1][2]  (.D(\input_filter[4][1] [2]), .CK(n_53_6), 
      .Q(\buffer[6][4][1] [2]), .QN());
   DFF_X1 \buffer_reg[6][4][1][1]  (.D(\input_filter[4][1] [1]), .CK(n_53_6), 
      .Q(\buffer[6][4][1] [1]), .QN());
   DFF_X1 \buffer_reg[6][4][1][0]  (.D(\input_filter[4][1] [0]), .CK(n_53_6), 
      .Q(\buffer[6][4][1] [0]), .QN());
   DFF_X1 \buffer_reg[5][4][1][15]  (.D(\input_filter[4][1] [15]), .CK(n_53_5), 
      .Q(\buffer[5][4][1] [15]), .QN());
   DFF_X1 \buffer_reg[5][4][1][14]  (.D(\input_filter[4][1] [14]), .CK(n_53_5), 
      .Q(\buffer[5][4][1] [14]), .QN());
   DFF_X1 \buffer_reg[5][4][1][13]  (.D(\input_filter[4][1] [13]), .CK(n_53_5), 
      .Q(\buffer[5][4][1] [13]), .QN());
   DFF_X1 \buffer_reg[5][4][1][12]  (.D(\input_filter[4][1] [12]), .CK(n_53_5), 
      .Q(\buffer[5][4][1] [12]), .QN());
   DFF_X1 \buffer_reg[5][4][1][11]  (.D(\input_filter[4][1] [11]), .CK(n_53_5), 
      .Q(\buffer[5][4][1] [11]), .QN());
   DFF_X1 \buffer_reg[5][4][1][10]  (.D(\input_filter[4][1] [10]), .CK(n_53_5), 
      .Q(\buffer[5][4][1] [10]), .QN());
   DFF_X1 \buffer_reg[5][4][1][9]  (.D(\input_filter[4][1] [9]), .CK(n_53_5), 
      .Q(\buffer[5][4][1] [9]), .QN());
   DFF_X1 \buffer_reg[5][4][1][8]  (.D(\input_filter[4][1] [8]), .CK(n_53_5), 
      .Q(\buffer[5][4][1] [8]), .QN());
   DFF_X1 \buffer_reg[5][4][1][7]  (.D(\input_filter[4][1] [7]), .CK(n_53_5), 
      .Q(\buffer[5][4][1] [7]), .QN());
   DFF_X1 \buffer_reg[5][4][1][6]  (.D(\input_filter[4][1] [6]), .CK(n_53_5), 
      .Q(\buffer[5][4][1] [6]), .QN());
   DFF_X1 \buffer_reg[5][4][1][5]  (.D(\input_filter[4][1] [5]), .CK(n_53_5), 
      .Q(\buffer[5][4][1] [5]), .QN());
   DFF_X1 \buffer_reg[5][4][1][4]  (.D(\input_filter[4][1] [4]), .CK(n_53_5), 
      .Q(\buffer[5][4][1] [4]), .QN());
   DFF_X1 \buffer_reg[5][4][1][3]  (.D(\input_filter[4][1] [3]), .CK(n_53_5), 
      .Q(\buffer[5][4][1] [3]), .QN());
   DFF_X1 \buffer_reg[5][4][1][2]  (.D(\input_filter[4][1] [2]), .CK(n_53_5), 
      .Q(\buffer[5][4][1] [2]), .QN());
   DFF_X1 \buffer_reg[5][4][1][1]  (.D(\input_filter[4][1] [1]), .CK(n_53_5), 
      .Q(\buffer[5][4][1] [1]), .QN());
   DFF_X1 \buffer_reg[5][4][1][0]  (.D(\input_filter[4][1] [0]), .CK(n_53_5), 
      .Q(\buffer[5][4][1] [0]), .QN());
   DFF_X1 \buffer_reg[4][4][1][15]  (.D(\input_filter[4][1] [15]), .CK(n_53_4), 
      .Q(\buffer[4][4][1] [15]), .QN());
   DFF_X1 \buffer_reg[4][4][1][14]  (.D(\input_filter[4][1] [14]), .CK(n_53_4), 
      .Q(\buffer[4][4][1] [14]), .QN());
   DFF_X1 \buffer_reg[4][4][1][13]  (.D(\input_filter[4][1] [13]), .CK(n_53_4), 
      .Q(\buffer[4][4][1] [13]), .QN());
   DFF_X1 \buffer_reg[4][4][1][12]  (.D(\input_filter[4][1] [12]), .CK(n_53_4), 
      .Q(\buffer[4][4][1] [12]), .QN());
   DFF_X1 \buffer_reg[4][4][1][11]  (.D(\input_filter[4][1] [11]), .CK(n_53_4), 
      .Q(\buffer[4][4][1] [11]), .QN());
   DFF_X1 \buffer_reg[4][4][1][10]  (.D(\input_filter[4][1] [10]), .CK(n_53_4), 
      .Q(\buffer[4][4][1] [10]), .QN());
   DFF_X1 \buffer_reg[4][4][1][9]  (.D(\input_filter[4][1] [9]), .CK(n_53_4), 
      .Q(\buffer[4][4][1] [9]), .QN());
   DFF_X1 \buffer_reg[4][4][1][8]  (.D(\input_filter[4][1] [8]), .CK(n_53_4), 
      .Q(\buffer[4][4][1] [8]), .QN());
   DFF_X1 \buffer_reg[4][4][1][7]  (.D(\input_filter[4][1] [7]), .CK(n_53_4), 
      .Q(\buffer[4][4][1] [7]), .QN());
   DFF_X1 \buffer_reg[4][4][1][6]  (.D(\input_filter[4][1] [6]), .CK(n_53_4), 
      .Q(\buffer[4][4][1] [6]), .QN());
   DFF_X1 \buffer_reg[4][4][1][5]  (.D(\input_filter[4][1] [5]), .CK(n_53_4), 
      .Q(\buffer[4][4][1] [5]), .QN());
   DFF_X1 \buffer_reg[4][4][1][4]  (.D(\input_filter[4][1] [4]), .CK(n_53_4), 
      .Q(\buffer[4][4][1] [4]), .QN());
   DFF_X1 \buffer_reg[4][4][1][3]  (.D(\input_filter[4][1] [3]), .CK(n_53_4), 
      .Q(\buffer[4][4][1] [3]), .QN());
   DFF_X1 \buffer_reg[4][4][1][2]  (.D(\input_filter[4][1] [2]), .CK(n_53_4), 
      .Q(\buffer[4][4][1] [2]), .QN());
   DFF_X1 \buffer_reg[4][4][1][1]  (.D(\input_filter[4][1] [1]), .CK(n_53_4), 
      .Q(\buffer[4][4][1] [1]), .QN());
   DFF_X1 \buffer_reg[4][4][1][0]  (.D(\input_filter[4][1] [0]), .CK(n_53_4), 
      .Q(\buffer[4][4][1] [0]), .QN());
   DFF_X1 \buffer_reg[3][4][1][15]  (.D(\input_filter[4][1] [15]), .CK(n_53_3), 
      .Q(\buffer[3][4][1] [15]), .QN());
   DFF_X1 \buffer_reg[3][4][1][14]  (.D(\input_filter[4][1] [14]), .CK(n_53_3), 
      .Q(\buffer[3][4][1] [14]), .QN());
   DFF_X1 \buffer_reg[3][4][1][13]  (.D(\input_filter[4][1] [13]), .CK(n_53_3), 
      .Q(\buffer[3][4][1] [13]), .QN());
   DFF_X1 \buffer_reg[3][4][1][12]  (.D(\input_filter[4][1] [12]), .CK(n_53_3), 
      .Q(\buffer[3][4][1] [12]), .QN());
   DFF_X1 \buffer_reg[3][4][1][11]  (.D(\input_filter[4][1] [11]), .CK(n_53_3), 
      .Q(\buffer[3][4][1] [11]), .QN());
   DFF_X1 \buffer_reg[3][4][1][10]  (.D(\input_filter[4][1] [10]), .CK(n_53_3), 
      .Q(\buffer[3][4][1] [10]), .QN());
   DFF_X1 \buffer_reg[3][4][1][9]  (.D(\input_filter[4][1] [9]), .CK(n_53_3), 
      .Q(\buffer[3][4][1] [9]), .QN());
   DFF_X1 \buffer_reg[3][4][1][8]  (.D(\input_filter[4][1] [8]), .CK(n_53_3), 
      .Q(\buffer[3][4][1] [8]), .QN());
   DFF_X1 \buffer_reg[3][4][1][7]  (.D(\input_filter[4][1] [7]), .CK(n_53_3), 
      .Q(\buffer[3][4][1] [7]), .QN());
   DFF_X1 \buffer_reg[3][4][1][6]  (.D(\input_filter[4][1] [6]), .CK(n_53_3), 
      .Q(\buffer[3][4][1] [6]), .QN());
   DFF_X1 \buffer_reg[3][4][1][5]  (.D(\input_filter[4][1] [5]), .CK(n_53_3), 
      .Q(\buffer[3][4][1] [5]), .QN());
   DFF_X1 \buffer_reg[3][4][1][4]  (.D(\input_filter[4][1] [4]), .CK(n_53_3), 
      .Q(\buffer[3][4][1] [4]), .QN());
   DFF_X1 \buffer_reg[3][4][1][3]  (.D(\input_filter[4][1] [3]), .CK(n_53_3), 
      .Q(\buffer[3][4][1] [3]), .QN());
   DFF_X1 \buffer_reg[3][4][1][2]  (.D(\input_filter[4][1] [2]), .CK(n_53_3), 
      .Q(\buffer[3][4][1] [2]), .QN());
   DFF_X1 \buffer_reg[3][4][1][1]  (.D(\input_filter[4][1] [1]), .CK(n_53_3), 
      .Q(\buffer[3][4][1] [1]), .QN());
   DFF_X1 \buffer_reg[3][4][1][0]  (.D(\input_filter[4][1] [0]), .CK(n_53_3), 
      .Q(\buffer[3][4][1] [0]), .QN());
   DFF_X1 \buffer_reg[2][4][1][15]  (.D(\input_filter[4][1] [15]), .CK(n_53_2), 
      .Q(\buffer[2][4][1] [15]), .QN());
   DFF_X1 \buffer_reg[2][4][1][14]  (.D(\input_filter[4][1] [14]), .CK(n_53_2), 
      .Q(\buffer[2][4][1] [14]), .QN());
   DFF_X1 \buffer_reg[2][4][1][13]  (.D(\input_filter[4][1] [13]), .CK(n_53_2), 
      .Q(\buffer[2][4][1] [13]), .QN());
   DFF_X1 \buffer_reg[2][4][1][12]  (.D(\input_filter[4][1] [12]), .CK(n_53_2), 
      .Q(\buffer[2][4][1] [12]), .QN());
   DFF_X1 \buffer_reg[2][4][1][11]  (.D(\input_filter[4][1] [11]), .CK(n_53_2), 
      .Q(\buffer[2][4][1] [11]), .QN());
   DFF_X1 \buffer_reg[2][4][1][10]  (.D(\input_filter[4][1] [10]), .CK(n_53_2), 
      .Q(\buffer[2][4][1] [10]), .QN());
   DFF_X1 \buffer_reg[2][4][1][9]  (.D(\input_filter[4][1] [9]), .CK(n_53_2), 
      .Q(\buffer[2][4][1] [9]), .QN());
   DFF_X1 \buffer_reg[2][4][1][8]  (.D(\input_filter[4][1] [8]), .CK(n_53_2), 
      .Q(\buffer[2][4][1] [8]), .QN());
   DFF_X1 \buffer_reg[2][4][1][7]  (.D(\input_filter[4][1] [7]), .CK(n_53_2), 
      .Q(\buffer[2][4][1] [7]), .QN());
   DFF_X1 \buffer_reg[2][4][1][6]  (.D(\input_filter[4][1] [6]), .CK(n_53_2), 
      .Q(\buffer[2][4][1] [6]), .QN());
   DFF_X1 \buffer_reg[2][4][1][5]  (.D(\input_filter[4][1] [5]), .CK(n_53_2), 
      .Q(\buffer[2][4][1] [5]), .QN());
   DFF_X1 \buffer_reg[2][4][1][4]  (.D(\input_filter[4][1] [4]), .CK(n_53_2), 
      .Q(\buffer[2][4][1] [4]), .QN());
   DFF_X1 \buffer_reg[2][4][1][3]  (.D(\input_filter[4][1] [3]), .CK(n_53_2), 
      .Q(\buffer[2][4][1] [3]), .QN());
   DFF_X1 \buffer_reg[2][4][1][2]  (.D(\input_filter[4][1] [2]), .CK(n_53_2), 
      .Q(\buffer[2][4][1] [2]), .QN());
   DFF_X1 \buffer_reg[2][4][1][1]  (.D(\input_filter[4][1] [1]), .CK(n_53_2), 
      .Q(\buffer[2][4][1] [1]), .QN());
   DFF_X1 \buffer_reg[2][4][1][0]  (.D(\input_filter[4][1] [0]), .CK(n_53_2), 
      .Q(\buffer[2][4][1] [0]), .QN());
   DFF_X1 \buffer_reg[1][4][1][15]  (.D(\input_filter[4][1] [15]), .CK(n_53_1), 
      .Q(\buffer[1][4][1] [15]), .QN());
   DFF_X1 \buffer_reg[1][4][1][14]  (.D(\input_filter[4][1] [14]), .CK(n_53_1), 
      .Q(\buffer[1][4][1] [14]), .QN());
   DFF_X1 \buffer_reg[1][4][1][13]  (.D(\input_filter[4][1] [13]), .CK(n_53_1), 
      .Q(\buffer[1][4][1] [13]), .QN());
   DFF_X1 \buffer_reg[1][4][1][12]  (.D(\input_filter[4][1] [12]), .CK(n_53_1), 
      .Q(\buffer[1][4][1] [12]), .QN());
   DFF_X1 \buffer_reg[1][4][1][11]  (.D(\input_filter[4][1] [11]), .CK(n_53_1), 
      .Q(\buffer[1][4][1] [11]), .QN());
   DFF_X1 \buffer_reg[1][4][1][10]  (.D(\input_filter[4][1] [10]), .CK(n_53_1), 
      .Q(\buffer[1][4][1] [10]), .QN());
   DFF_X1 \buffer_reg[1][4][1][9]  (.D(\input_filter[4][1] [9]), .CK(n_53_1), 
      .Q(\buffer[1][4][1] [9]), .QN());
   DFF_X1 \buffer_reg[1][4][1][8]  (.D(\input_filter[4][1] [8]), .CK(n_53_1), 
      .Q(\buffer[1][4][1] [8]), .QN());
   DFF_X1 \buffer_reg[1][4][1][7]  (.D(\input_filter[4][1] [7]), .CK(n_53_1), 
      .Q(\buffer[1][4][1] [7]), .QN());
   DFF_X1 \buffer_reg[1][4][1][6]  (.D(\input_filter[4][1] [6]), .CK(n_53_1), 
      .Q(\buffer[1][4][1] [6]), .QN());
   DFF_X1 \buffer_reg[1][4][1][5]  (.D(\input_filter[4][1] [5]), .CK(n_53_1), 
      .Q(\buffer[1][4][1] [5]), .QN());
   DFF_X1 \buffer_reg[1][4][1][4]  (.D(\input_filter[4][1] [4]), .CK(n_53_1), 
      .Q(\buffer[1][4][1] [4]), .QN());
   DFF_X1 \buffer_reg[1][4][1][3]  (.D(\input_filter[4][1] [3]), .CK(n_53_1), 
      .Q(\buffer[1][4][1] [3]), .QN());
   DFF_X1 \buffer_reg[1][4][1][2]  (.D(\input_filter[4][1] [2]), .CK(n_53_1), 
      .Q(\buffer[1][4][1] [2]), .QN());
   DFF_X1 \buffer_reg[1][4][1][1]  (.D(\input_filter[4][1] [1]), .CK(n_53_1), 
      .Q(\buffer[1][4][1] [1]), .QN());
   DFF_X1 \buffer_reg[1][4][1][0]  (.D(\input_filter[4][1] [0]), .CK(n_53_1), 
      .Q(\buffer[1][4][1] [0]), .QN());
   DFF_X1 \buffer_reg[0][4][1][15]  (.D(\input_filter[4][1] [15]), .CK(n_53_0), 
      .Q(\buffer[0][4][1] [15]), .QN());
   DFF_X1 \buffer_reg[0][4][1][14]  (.D(\input_filter[4][1] [14]), .CK(n_53_0), 
      .Q(\buffer[0][4][1] [14]), .QN());
   DFF_X1 \buffer_reg[0][4][1][13]  (.D(\input_filter[4][1] [13]), .CK(n_53_0), 
      .Q(\buffer[0][4][1] [13]), .QN());
   DFF_X1 \buffer_reg[0][4][1][12]  (.D(\input_filter[4][1] [12]), .CK(n_53_0), 
      .Q(\buffer[0][4][1] [12]), .QN());
   DFF_X1 \buffer_reg[0][4][1][11]  (.D(\input_filter[4][1] [11]), .CK(n_53_0), 
      .Q(\buffer[0][4][1] [11]), .QN());
   DFF_X1 \buffer_reg[0][4][1][10]  (.D(\input_filter[4][1] [10]), .CK(n_53_0), 
      .Q(\buffer[0][4][1] [10]), .QN());
   DFF_X1 \buffer_reg[0][4][1][9]  (.D(\input_filter[4][1] [9]), .CK(n_53_0), 
      .Q(\buffer[0][4][1] [9]), .QN());
   DFF_X1 \buffer_reg[0][4][1][8]  (.D(\input_filter[4][1] [8]), .CK(n_53_0), 
      .Q(\buffer[0][4][1] [8]), .QN());
   DFF_X1 \buffer_reg[0][4][1][7]  (.D(\input_filter[4][1] [7]), .CK(n_53_0), 
      .Q(\buffer[0][4][1] [7]), .QN());
   DFF_X1 \buffer_reg[0][4][1][6]  (.D(\input_filter[4][1] [6]), .CK(n_53_0), 
      .Q(\buffer[0][4][1] [6]), .QN());
   DFF_X1 \buffer_reg[0][4][1][5]  (.D(\input_filter[4][1] [5]), .CK(n_53_0), 
      .Q(\buffer[0][4][1] [5]), .QN());
   DFF_X1 \buffer_reg[0][4][1][4]  (.D(\input_filter[4][1] [4]), .CK(n_53_0), 
      .Q(\buffer[0][4][1] [4]), .QN());
   DFF_X1 \buffer_reg[0][4][1][3]  (.D(\input_filter[4][1] [3]), .CK(n_53_0), 
      .Q(\buffer[0][4][1] [3]), .QN());
   DFF_X1 \buffer_reg[0][4][1][2]  (.D(\input_filter[4][1] [2]), .CK(n_53_0), 
      .Q(\buffer[0][4][1] [2]), .QN());
   DFF_X1 \buffer_reg[0][4][1][1]  (.D(\input_filter[4][1] [1]), .CK(n_53_0), 
      .Q(\buffer[0][4][1] [1]), .QN());
   DFF_X1 \buffer_reg[0][4][1][0]  (.D(\input_filter[4][1] [0]), .CK(n_53_0), 
      .Q(\buffer[0][4][1] [0]), .QN());
   DFF_X1 \buffer_reg[15][4][0][15]  (.D(\input_filter[4][0] [15]), .CK(n_53_15), 
      .Q(\buffer[15][4][0] [15]), .QN());
   DFF_X1 \buffer_reg[15][4][0][14]  (.D(\input_filter[4][0] [14]), .CK(n_53_15), 
      .Q(\buffer[15][4][0] [14]), .QN());
   DFF_X1 \buffer_reg[15][4][0][13]  (.D(\input_filter[4][0] [13]), .CK(n_53_15), 
      .Q(\buffer[15][4][0] [13]), .QN());
   DFF_X1 \buffer_reg[15][4][0][12]  (.D(\input_filter[4][0] [12]), .CK(n_53_15), 
      .Q(\buffer[15][4][0] [12]), .QN());
   DFF_X1 \buffer_reg[15][4][0][11]  (.D(\input_filter[4][0] [11]), .CK(n_53_15), 
      .Q(\buffer[15][4][0] [11]), .QN());
   DFF_X1 \buffer_reg[15][4][0][10]  (.D(\input_filter[4][0] [10]), .CK(n_53_15), 
      .Q(\buffer[15][4][0] [10]), .QN());
   DFF_X1 \buffer_reg[15][4][0][9]  (.D(\input_filter[4][0] [9]), .CK(n_53_15), 
      .Q(\buffer[15][4][0] [9]), .QN());
   DFF_X1 \buffer_reg[15][4][0][8]  (.D(\input_filter[4][0] [8]), .CK(n_53_15), 
      .Q(\buffer[15][4][0] [8]), .QN());
   DFF_X1 \buffer_reg[15][4][0][7]  (.D(\input_filter[4][0] [7]), .CK(n_53_15), 
      .Q(\buffer[15][4][0] [7]), .QN());
   DFF_X1 \buffer_reg[15][4][0][6]  (.D(\input_filter[4][0] [6]), .CK(n_53_15), 
      .Q(\buffer[15][4][0] [6]), .QN());
   DFF_X1 \buffer_reg[15][4][0][5]  (.D(\input_filter[4][0] [5]), .CK(n_53_15), 
      .Q(\buffer[15][4][0] [5]), .QN());
   DFF_X1 \buffer_reg[15][4][0][4]  (.D(\input_filter[4][0] [4]), .CK(n_53_15), 
      .Q(\buffer[15][4][0] [4]), .QN());
   DFF_X1 \buffer_reg[15][4][0][3]  (.D(\input_filter[4][0] [3]), .CK(n_53_15), 
      .Q(\buffer[15][4][0] [3]), .QN());
   DFF_X1 \buffer_reg[15][4][0][2]  (.D(\input_filter[4][0] [2]), .CK(n_53_15), 
      .Q(\buffer[15][4][0] [2]), .QN());
   DFF_X1 \buffer_reg[15][4][0][1]  (.D(\input_filter[4][0] [1]), .CK(n_53_15), 
      .Q(\buffer[15][4][0] [1]), .QN());
   DFF_X1 \buffer_reg[15][4][0][0]  (.D(\input_filter[4][0] [0]), .CK(n_53_15), 
      .Q(\buffer[15][4][0] [0]), .QN());
   DFF_X1 \buffer_reg[14][4][0][15]  (.D(\input_filter[4][0] [15]), .CK(n_53_14), 
      .Q(\buffer[14][4][0] [15]), .QN());
   DFF_X1 \buffer_reg[14][4][0][14]  (.D(\input_filter[4][0] [14]), .CK(n_53_14), 
      .Q(\buffer[14][4][0] [14]), .QN());
   DFF_X1 \buffer_reg[14][4][0][13]  (.D(\input_filter[4][0] [13]), .CK(n_53_14), 
      .Q(\buffer[14][4][0] [13]), .QN());
   DFF_X1 \buffer_reg[14][4][0][12]  (.D(\input_filter[4][0] [12]), .CK(n_53_14), 
      .Q(\buffer[14][4][0] [12]), .QN());
   DFF_X1 \buffer_reg[14][4][0][11]  (.D(\input_filter[4][0] [11]), .CK(n_53_14), 
      .Q(\buffer[14][4][0] [11]), .QN());
   DFF_X1 \buffer_reg[14][4][0][10]  (.D(\input_filter[4][0] [10]), .CK(n_53_14), 
      .Q(\buffer[14][4][0] [10]), .QN());
   DFF_X1 \buffer_reg[14][4][0][9]  (.D(\input_filter[4][0] [9]), .CK(n_53_14), 
      .Q(\buffer[14][4][0] [9]), .QN());
   DFF_X1 \buffer_reg[14][4][0][8]  (.D(\input_filter[4][0] [8]), .CK(n_53_14), 
      .Q(\buffer[14][4][0] [8]), .QN());
   DFF_X1 \buffer_reg[14][4][0][7]  (.D(\input_filter[4][0] [7]), .CK(n_53_14), 
      .Q(\buffer[14][4][0] [7]), .QN());
   DFF_X1 \buffer_reg[14][4][0][6]  (.D(\input_filter[4][0] [6]), .CK(n_53_14), 
      .Q(\buffer[14][4][0] [6]), .QN());
   DFF_X1 \buffer_reg[14][4][0][5]  (.D(\input_filter[4][0] [5]), .CK(n_53_14), 
      .Q(\buffer[14][4][0] [5]), .QN());
   DFF_X1 \buffer_reg[14][4][0][4]  (.D(\input_filter[4][0] [4]), .CK(n_53_14), 
      .Q(\buffer[14][4][0] [4]), .QN());
   DFF_X1 \buffer_reg[14][4][0][3]  (.D(\input_filter[4][0] [3]), .CK(n_53_14), 
      .Q(\buffer[14][4][0] [3]), .QN());
   DFF_X1 \buffer_reg[14][4][0][2]  (.D(\input_filter[4][0] [2]), .CK(n_53_14), 
      .Q(\buffer[14][4][0] [2]), .QN());
   DFF_X1 \buffer_reg[14][4][0][1]  (.D(\input_filter[4][0] [1]), .CK(n_53_14), 
      .Q(\buffer[14][4][0] [1]), .QN());
   DFF_X1 \buffer_reg[14][4][0][0]  (.D(\input_filter[4][0] [0]), .CK(n_53_14), 
      .Q(\buffer[14][4][0] [0]), .QN());
   DFF_X1 \buffer_reg[13][4][0][15]  (.D(\input_filter[4][0] [15]), .CK(n_53_13), 
      .Q(\buffer[13][4][0] [15]), .QN());
   DFF_X1 \buffer_reg[13][4][0][14]  (.D(\input_filter[4][0] [14]), .CK(n_53_13), 
      .Q(\buffer[13][4][0] [14]), .QN());
   DFF_X1 \buffer_reg[13][4][0][13]  (.D(\input_filter[4][0] [13]), .CK(n_53_13), 
      .Q(\buffer[13][4][0] [13]), .QN());
   DFF_X1 \buffer_reg[13][4][0][12]  (.D(\input_filter[4][0] [12]), .CK(n_53_13), 
      .Q(\buffer[13][4][0] [12]), .QN());
   DFF_X1 \buffer_reg[13][4][0][11]  (.D(\input_filter[4][0] [11]), .CK(n_53_13), 
      .Q(\buffer[13][4][0] [11]), .QN());
   DFF_X1 \buffer_reg[13][4][0][10]  (.D(\input_filter[4][0] [10]), .CK(n_53_13), 
      .Q(\buffer[13][4][0] [10]), .QN());
   DFF_X1 \buffer_reg[13][4][0][9]  (.D(\input_filter[4][0] [9]), .CK(n_53_13), 
      .Q(\buffer[13][4][0] [9]), .QN());
   DFF_X1 \buffer_reg[13][4][0][8]  (.D(\input_filter[4][0] [8]), .CK(n_53_13), 
      .Q(\buffer[13][4][0] [8]), .QN());
   DFF_X1 \buffer_reg[13][4][0][7]  (.D(\input_filter[4][0] [7]), .CK(n_53_13), 
      .Q(\buffer[13][4][0] [7]), .QN());
   DFF_X1 \buffer_reg[13][4][0][6]  (.D(\input_filter[4][0] [6]), .CK(n_53_13), 
      .Q(\buffer[13][4][0] [6]), .QN());
   DFF_X1 \buffer_reg[13][4][0][5]  (.D(\input_filter[4][0] [5]), .CK(n_53_13), 
      .Q(\buffer[13][4][0] [5]), .QN());
   DFF_X1 \buffer_reg[13][4][0][4]  (.D(\input_filter[4][0] [4]), .CK(n_53_13), 
      .Q(\buffer[13][4][0] [4]), .QN());
   DFF_X1 \buffer_reg[13][4][0][3]  (.D(\input_filter[4][0] [3]), .CK(n_53_13), 
      .Q(\buffer[13][4][0] [3]), .QN());
   DFF_X1 \buffer_reg[13][4][0][2]  (.D(\input_filter[4][0] [2]), .CK(n_53_13), 
      .Q(\buffer[13][4][0] [2]), .QN());
   DFF_X1 \buffer_reg[13][4][0][1]  (.D(\input_filter[4][0] [1]), .CK(n_53_13), 
      .Q(\buffer[13][4][0] [1]), .QN());
   DFF_X1 \buffer_reg[13][4][0][0]  (.D(\input_filter[4][0] [0]), .CK(n_53_13), 
      .Q(\buffer[13][4][0] [0]), .QN());
   DFF_X1 \buffer_reg[12][4][0][15]  (.D(\input_filter[4][0] [15]), .CK(n_53_12), 
      .Q(\buffer[12][4][0] [15]), .QN());
   DFF_X1 \buffer_reg[12][4][0][14]  (.D(\input_filter[4][0] [14]), .CK(n_53_12), 
      .Q(\buffer[12][4][0] [14]), .QN());
   DFF_X1 \buffer_reg[12][4][0][13]  (.D(\input_filter[4][0] [13]), .CK(n_53_12), 
      .Q(\buffer[12][4][0] [13]), .QN());
   DFF_X1 \buffer_reg[12][4][0][12]  (.D(\input_filter[4][0] [12]), .CK(n_53_12), 
      .Q(\buffer[12][4][0] [12]), .QN());
   DFF_X1 \buffer_reg[12][4][0][11]  (.D(\input_filter[4][0] [11]), .CK(n_53_12), 
      .Q(\buffer[12][4][0] [11]), .QN());
   DFF_X1 \buffer_reg[12][4][0][10]  (.D(\input_filter[4][0] [10]), .CK(n_53_12), 
      .Q(\buffer[12][4][0] [10]), .QN());
   DFF_X1 \buffer_reg[12][4][0][9]  (.D(\input_filter[4][0] [9]), .CK(n_53_12), 
      .Q(\buffer[12][4][0] [9]), .QN());
   DFF_X1 \buffer_reg[12][4][0][8]  (.D(\input_filter[4][0] [8]), .CK(n_53_12), 
      .Q(\buffer[12][4][0] [8]), .QN());
   DFF_X1 \buffer_reg[12][4][0][7]  (.D(\input_filter[4][0] [7]), .CK(n_53_12), 
      .Q(\buffer[12][4][0] [7]), .QN());
   DFF_X1 \buffer_reg[12][4][0][6]  (.D(\input_filter[4][0] [6]), .CK(n_53_12), 
      .Q(\buffer[12][4][0] [6]), .QN());
   DFF_X1 \buffer_reg[12][4][0][5]  (.D(\input_filter[4][0] [5]), .CK(n_53_12), 
      .Q(\buffer[12][4][0] [5]), .QN());
   DFF_X1 \buffer_reg[12][4][0][4]  (.D(\input_filter[4][0] [4]), .CK(n_53_12), 
      .Q(\buffer[12][4][0] [4]), .QN());
   DFF_X1 \buffer_reg[12][4][0][3]  (.D(\input_filter[4][0] [3]), .CK(n_53_12), 
      .Q(\buffer[12][4][0] [3]), .QN());
   DFF_X1 \buffer_reg[12][4][0][2]  (.D(\input_filter[4][0] [2]), .CK(n_53_12), 
      .Q(\buffer[12][4][0] [2]), .QN());
   DFF_X1 \buffer_reg[12][4][0][1]  (.D(\input_filter[4][0] [1]), .CK(n_53_12), 
      .Q(\buffer[12][4][0] [1]), .QN());
   DFF_X1 \buffer_reg[12][4][0][0]  (.D(\input_filter[4][0] [0]), .CK(n_53_12), 
      .Q(\buffer[12][4][0] [0]), .QN());
   DFF_X1 \buffer_reg[11][4][0][15]  (.D(\input_filter[4][0] [15]), .CK(n_53_11), 
      .Q(\buffer[11][4][0] [15]), .QN());
   DFF_X1 \buffer_reg[11][4][0][14]  (.D(\input_filter[4][0] [14]), .CK(n_53_11), 
      .Q(\buffer[11][4][0] [14]), .QN());
   DFF_X1 \buffer_reg[11][4][0][13]  (.D(\input_filter[4][0] [13]), .CK(n_53_11), 
      .Q(\buffer[11][4][0] [13]), .QN());
   DFF_X1 \buffer_reg[11][4][0][12]  (.D(\input_filter[4][0] [12]), .CK(n_53_11), 
      .Q(\buffer[11][4][0] [12]), .QN());
   DFF_X1 \buffer_reg[11][4][0][11]  (.D(\input_filter[4][0] [11]), .CK(n_53_11), 
      .Q(\buffer[11][4][0] [11]), .QN());
   DFF_X1 \buffer_reg[11][4][0][10]  (.D(\input_filter[4][0] [10]), .CK(n_53_11), 
      .Q(\buffer[11][4][0] [10]), .QN());
   DFF_X1 \buffer_reg[11][4][0][9]  (.D(\input_filter[4][0] [9]), .CK(n_53_11), 
      .Q(\buffer[11][4][0] [9]), .QN());
   DFF_X1 \buffer_reg[11][4][0][8]  (.D(\input_filter[4][0] [8]), .CK(n_53_11), 
      .Q(\buffer[11][4][0] [8]), .QN());
   DFF_X1 \buffer_reg[11][4][0][7]  (.D(\input_filter[4][0] [7]), .CK(n_53_11), 
      .Q(\buffer[11][4][0] [7]), .QN());
   DFF_X1 \buffer_reg[11][4][0][6]  (.D(\input_filter[4][0] [6]), .CK(n_53_11), 
      .Q(\buffer[11][4][0] [6]), .QN());
   DFF_X1 \buffer_reg[11][4][0][5]  (.D(\input_filter[4][0] [5]), .CK(n_53_11), 
      .Q(\buffer[11][4][0] [5]), .QN());
   DFF_X1 \buffer_reg[11][4][0][4]  (.D(\input_filter[4][0] [4]), .CK(n_53_11), 
      .Q(\buffer[11][4][0] [4]), .QN());
   DFF_X1 \buffer_reg[11][4][0][3]  (.D(\input_filter[4][0] [3]), .CK(n_53_11), 
      .Q(\buffer[11][4][0] [3]), .QN());
   DFF_X1 \buffer_reg[11][4][0][2]  (.D(\input_filter[4][0] [2]), .CK(n_53_11), 
      .Q(\buffer[11][4][0] [2]), .QN());
   DFF_X1 \buffer_reg[11][4][0][1]  (.D(\input_filter[4][0] [1]), .CK(n_53_11), 
      .Q(\buffer[11][4][0] [1]), .QN());
   DFF_X1 \buffer_reg[11][4][0][0]  (.D(\input_filter[4][0] [0]), .CK(n_53_11), 
      .Q(\buffer[11][4][0] [0]), .QN());
   DFF_X1 \buffer_reg[10][4][0][15]  (.D(\input_filter[4][0] [15]), .CK(n_53_10), 
      .Q(\buffer[10][4][0] [15]), .QN());
   DFF_X1 \buffer_reg[10][4][0][14]  (.D(\input_filter[4][0] [14]), .CK(n_53_10), 
      .Q(\buffer[10][4][0] [14]), .QN());
   DFF_X1 \buffer_reg[10][4][0][13]  (.D(\input_filter[4][0] [13]), .CK(n_53_10), 
      .Q(\buffer[10][4][0] [13]), .QN());
   DFF_X1 \buffer_reg[10][4][0][12]  (.D(\input_filter[4][0] [12]), .CK(n_53_10), 
      .Q(\buffer[10][4][0] [12]), .QN());
   DFF_X1 \buffer_reg[10][4][0][11]  (.D(\input_filter[4][0] [11]), .CK(n_53_10), 
      .Q(\buffer[10][4][0] [11]), .QN());
   DFF_X1 \buffer_reg[10][4][0][10]  (.D(\input_filter[4][0] [10]), .CK(n_53_10), 
      .Q(\buffer[10][4][0] [10]), .QN());
   DFF_X1 \buffer_reg[10][4][0][9]  (.D(\input_filter[4][0] [9]), .CK(n_53_10), 
      .Q(\buffer[10][4][0] [9]), .QN());
   DFF_X1 \buffer_reg[10][4][0][8]  (.D(\input_filter[4][0] [8]), .CK(n_53_10), 
      .Q(\buffer[10][4][0] [8]), .QN());
   DFF_X1 \buffer_reg[10][4][0][7]  (.D(\input_filter[4][0] [7]), .CK(n_53_10), 
      .Q(\buffer[10][4][0] [7]), .QN());
   DFF_X1 \buffer_reg[10][4][0][6]  (.D(\input_filter[4][0] [6]), .CK(n_53_10), 
      .Q(\buffer[10][4][0] [6]), .QN());
   DFF_X1 \buffer_reg[10][4][0][5]  (.D(\input_filter[4][0] [5]), .CK(n_53_10), 
      .Q(\buffer[10][4][0] [5]), .QN());
   DFF_X1 \buffer_reg[10][4][0][4]  (.D(\input_filter[4][0] [4]), .CK(n_53_10), 
      .Q(\buffer[10][4][0] [4]), .QN());
   DFF_X1 \buffer_reg[10][4][0][3]  (.D(\input_filter[4][0] [3]), .CK(n_53_10), 
      .Q(\buffer[10][4][0] [3]), .QN());
   DFF_X1 \buffer_reg[10][4][0][2]  (.D(\input_filter[4][0] [2]), .CK(n_53_10), 
      .Q(\buffer[10][4][0] [2]), .QN());
   DFF_X1 \buffer_reg[10][4][0][1]  (.D(\input_filter[4][0] [1]), .CK(n_53_10), 
      .Q(\buffer[10][4][0] [1]), .QN());
   DFF_X1 \buffer_reg[10][4][0][0]  (.D(\input_filter[4][0] [0]), .CK(n_53_10), 
      .Q(\buffer[10][4][0] [0]), .QN());
   DFF_X1 \buffer_reg[9][4][0][15]  (.D(\input_filter[4][0] [15]), .CK(n_53_9), 
      .Q(\buffer[9][4][0] [15]), .QN());
   DFF_X1 \buffer_reg[9][4][0][14]  (.D(\input_filter[4][0] [14]), .CK(n_53_9), 
      .Q(\buffer[9][4][0] [14]), .QN());
   DFF_X1 \buffer_reg[9][4][0][13]  (.D(\input_filter[4][0] [13]), .CK(n_53_9), 
      .Q(\buffer[9][4][0] [13]), .QN());
   DFF_X1 \buffer_reg[9][4][0][12]  (.D(\input_filter[4][0] [12]), .CK(n_53_9), 
      .Q(\buffer[9][4][0] [12]), .QN());
   DFF_X1 \buffer_reg[9][4][0][11]  (.D(\input_filter[4][0] [11]), .CK(n_53_9), 
      .Q(\buffer[9][4][0] [11]), .QN());
   DFF_X1 \buffer_reg[9][4][0][10]  (.D(\input_filter[4][0] [10]), .CK(n_53_9), 
      .Q(\buffer[9][4][0] [10]), .QN());
   DFF_X1 \buffer_reg[9][4][0][9]  (.D(\input_filter[4][0] [9]), .CK(n_53_9), 
      .Q(\buffer[9][4][0] [9]), .QN());
   DFF_X1 \buffer_reg[9][4][0][8]  (.D(\input_filter[4][0] [8]), .CK(n_53_9), 
      .Q(\buffer[9][4][0] [8]), .QN());
   DFF_X1 \buffer_reg[9][4][0][7]  (.D(\input_filter[4][0] [7]), .CK(n_53_9), 
      .Q(\buffer[9][4][0] [7]), .QN());
   DFF_X1 \buffer_reg[9][4][0][6]  (.D(\input_filter[4][0] [6]), .CK(n_53_9), 
      .Q(\buffer[9][4][0] [6]), .QN());
   DFF_X1 \buffer_reg[9][4][0][5]  (.D(\input_filter[4][0] [5]), .CK(n_53_9), 
      .Q(\buffer[9][4][0] [5]), .QN());
   DFF_X1 \buffer_reg[9][4][0][4]  (.D(\input_filter[4][0] [4]), .CK(n_53_9), 
      .Q(\buffer[9][4][0] [4]), .QN());
   DFF_X1 \buffer_reg[9][4][0][3]  (.D(\input_filter[4][0] [3]), .CK(n_53_9), 
      .Q(\buffer[9][4][0] [3]), .QN());
   DFF_X1 \buffer_reg[9][4][0][2]  (.D(\input_filter[4][0] [2]), .CK(n_53_9), 
      .Q(\buffer[9][4][0] [2]), .QN());
   DFF_X1 \buffer_reg[9][4][0][1]  (.D(\input_filter[4][0] [1]), .CK(n_53_9), 
      .Q(\buffer[9][4][0] [1]), .QN());
   DFF_X1 \buffer_reg[9][4][0][0]  (.D(\input_filter[4][0] [0]), .CK(n_53_9), 
      .Q(\buffer[9][4][0] [0]), .QN());
   DFF_X1 \buffer_reg[8][4][0][15]  (.D(\input_filter[4][0] [15]), .CK(n_53_8), 
      .Q(\buffer[8][4][0] [15]), .QN());
   DFF_X1 \buffer_reg[8][4][0][14]  (.D(\input_filter[4][0] [14]), .CK(n_53_8), 
      .Q(\buffer[8][4][0] [14]), .QN());
   DFF_X1 \buffer_reg[8][4][0][13]  (.D(\input_filter[4][0] [13]), .CK(n_53_8), 
      .Q(\buffer[8][4][0] [13]), .QN());
   DFF_X1 \buffer_reg[8][4][0][12]  (.D(\input_filter[4][0] [12]), .CK(n_53_8), 
      .Q(\buffer[8][4][0] [12]), .QN());
   DFF_X1 \buffer_reg[8][4][0][11]  (.D(\input_filter[4][0] [11]), .CK(n_53_8), 
      .Q(\buffer[8][4][0] [11]), .QN());
   DFF_X1 \buffer_reg[8][4][0][10]  (.D(\input_filter[4][0] [10]), .CK(n_53_8), 
      .Q(\buffer[8][4][0] [10]), .QN());
   DFF_X1 \buffer_reg[8][4][0][9]  (.D(\input_filter[4][0] [9]), .CK(n_53_8), 
      .Q(\buffer[8][4][0] [9]), .QN());
   DFF_X1 \buffer_reg[8][4][0][8]  (.D(\input_filter[4][0] [8]), .CK(n_53_8), 
      .Q(\buffer[8][4][0] [8]), .QN());
   DFF_X1 \buffer_reg[8][4][0][7]  (.D(\input_filter[4][0] [7]), .CK(n_53_8), 
      .Q(\buffer[8][4][0] [7]), .QN());
   DFF_X1 \buffer_reg[8][4][0][6]  (.D(\input_filter[4][0] [6]), .CK(n_53_8), 
      .Q(\buffer[8][4][0] [6]), .QN());
   DFF_X1 \buffer_reg[8][4][0][5]  (.D(\input_filter[4][0] [5]), .CK(n_53_8), 
      .Q(\buffer[8][4][0] [5]), .QN());
   DFF_X1 \buffer_reg[8][4][0][4]  (.D(\input_filter[4][0] [4]), .CK(n_53_8), 
      .Q(\buffer[8][4][0] [4]), .QN());
   DFF_X1 \buffer_reg[8][4][0][3]  (.D(\input_filter[4][0] [3]), .CK(n_53_8), 
      .Q(\buffer[8][4][0] [3]), .QN());
   DFF_X1 \buffer_reg[8][4][0][2]  (.D(\input_filter[4][0] [2]), .CK(n_53_8), 
      .Q(\buffer[8][4][0] [2]), .QN());
   DFF_X1 \buffer_reg[8][4][0][1]  (.D(\input_filter[4][0] [1]), .CK(n_53_8), 
      .Q(\buffer[8][4][0] [1]), .QN());
   DFF_X1 \buffer_reg[8][4][0][0]  (.D(\input_filter[4][0] [0]), .CK(n_53_8), 
      .Q(\buffer[8][4][0] [0]), .QN());
   DFF_X1 \buffer_reg[7][4][0][15]  (.D(\input_filter[4][0] [15]), .CK(n_53_7), 
      .Q(\buffer[7][4][0] [15]), .QN());
   DFF_X1 \buffer_reg[7][4][0][14]  (.D(\input_filter[4][0] [14]), .CK(n_53_7), 
      .Q(\buffer[7][4][0] [14]), .QN());
   DFF_X1 \buffer_reg[7][4][0][13]  (.D(\input_filter[4][0] [13]), .CK(n_53_7), 
      .Q(\buffer[7][4][0] [13]), .QN());
   DFF_X1 \buffer_reg[7][4][0][12]  (.D(\input_filter[4][0] [12]), .CK(n_53_7), 
      .Q(\buffer[7][4][0] [12]), .QN());
   DFF_X1 \buffer_reg[7][4][0][11]  (.D(\input_filter[4][0] [11]), .CK(n_53_7), 
      .Q(\buffer[7][4][0] [11]), .QN());
   DFF_X1 \buffer_reg[7][4][0][10]  (.D(\input_filter[4][0] [10]), .CK(n_53_7), 
      .Q(\buffer[7][4][0] [10]), .QN());
   DFF_X1 \buffer_reg[7][4][0][9]  (.D(\input_filter[4][0] [9]), .CK(n_53_7), 
      .Q(\buffer[7][4][0] [9]), .QN());
   DFF_X1 \buffer_reg[7][4][0][8]  (.D(\input_filter[4][0] [8]), .CK(n_53_7), 
      .Q(\buffer[7][4][0] [8]), .QN());
   DFF_X1 \buffer_reg[7][4][0][7]  (.D(\input_filter[4][0] [7]), .CK(n_53_7), 
      .Q(\buffer[7][4][0] [7]), .QN());
   DFF_X1 \buffer_reg[7][4][0][6]  (.D(\input_filter[4][0] [6]), .CK(n_53_7), 
      .Q(\buffer[7][4][0] [6]), .QN());
   DFF_X1 \buffer_reg[7][4][0][5]  (.D(\input_filter[4][0] [5]), .CK(n_53_7), 
      .Q(\buffer[7][4][0] [5]), .QN());
   DFF_X1 \buffer_reg[7][4][0][4]  (.D(\input_filter[4][0] [4]), .CK(n_53_7), 
      .Q(\buffer[7][4][0] [4]), .QN());
   DFF_X1 \buffer_reg[7][4][0][3]  (.D(\input_filter[4][0] [3]), .CK(n_53_7), 
      .Q(\buffer[7][4][0] [3]), .QN());
   DFF_X1 \buffer_reg[7][4][0][2]  (.D(\input_filter[4][0] [2]), .CK(n_53_7), 
      .Q(\buffer[7][4][0] [2]), .QN());
   DFF_X1 \buffer_reg[7][4][0][1]  (.D(\input_filter[4][0] [1]), .CK(n_53_7), 
      .Q(\buffer[7][4][0] [1]), .QN());
   DFF_X1 \buffer_reg[7][4][0][0]  (.D(\input_filter[4][0] [0]), .CK(n_53_7), 
      .Q(\buffer[7][4][0] [0]), .QN());
   DFF_X1 \buffer_reg[6][4][0][15]  (.D(\input_filter[4][0] [15]), .CK(n_53_6), 
      .Q(\buffer[6][4][0] [15]), .QN());
   DFF_X1 \buffer_reg[6][4][0][14]  (.D(\input_filter[4][0] [14]), .CK(n_53_6), 
      .Q(\buffer[6][4][0] [14]), .QN());
   DFF_X1 \buffer_reg[6][4][0][13]  (.D(\input_filter[4][0] [13]), .CK(n_53_6), 
      .Q(\buffer[6][4][0] [13]), .QN());
   DFF_X1 \buffer_reg[6][4][0][12]  (.D(\input_filter[4][0] [12]), .CK(n_53_6), 
      .Q(\buffer[6][4][0] [12]), .QN());
   DFF_X1 \buffer_reg[6][4][0][11]  (.D(\input_filter[4][0] [11]), .CK(n_53_6), 
      .Q(\buffer[6][4][0] [11]), .QN());
   DFF_X1 \buffer_reg[6][4][0][10]  (.D(\input_filter[4][0] [10]), .CK(n_53_6), 
      .Q(\buffer[6][4][0] [10]), .QN());
   DFF_X1 \buffer_reg[6][4][0][9]  (.D(\input_filter[4][0] [9]), .CK(n_53_6), 
      .Q(\buffer[6][4][0] [9]), .QN());
   DFF_X1 \buffer_reg[6][4][0][8]  (.D(\input_filter[4][0] [8]), .CK(n_53_6), 
      .Q(\buffer[6][4][0] [8]), .QN());
   DFF_X1 \buffer_reg[6][4][0][7]  (.D(\input_filter[4][0] [7]), .CK(n_53_6), 
      .Q(\buffer[6][4][0] [7]), .QN());
   DFF_X1 \buffer_reg[6][4][0][6]  (.D(\input_filter[4][0] [6]), .CK(n_53_6), 
      .Q(\buffer[6][4][0] [6]), .QN());
   DFF_X1 \buffer_reg[6][4][0][5]  (.D(\input_filter[4][0] [5]), .CK(n_53_6), 
      .Q(\buffer[6][4][0] [5]), .QN());
   DFF_X1 \buffer_reg[6][4][0][4]  (.D(\input_filter[4][0] [4]), .CK(n_53_6), 
      .Q(\buffer[6][4][0] [4]), .QN());
   DFF_X1 \buffer_reg[6][4][0][3]  (.D(\input_filter[4][0] [3]), .CK(n_53_6), 
      .Q(\buffer[6][4][0] [3]), .QN());
   DFF_X1 \buffer_reg[6][4][0][2]  (.D(\input_filter[4][0] [2]), .CK(n_53_6), 
      .Q(\buffer[6][4][0] [2]), .QN());
   DFF_X1 \buffer_reg[6][4][0][1]  (.D(\input_filter[4][0] [1]), .CK(n_53_6), 
      .Q(\buffer[6][4][0] [1]), .QN());
   DFF_X1 \buffer_reg[6][4][0][0]  (.D(\input_filter[4][0] [0]), .CK(n_53_6), 
      .Q(\buffer[6][4][0] [0]), .QN());
   DFF_X1 \buffer_reg[5][4][0][15]  (.D(\input_filter[4][0] [15]), .CK(n_53_5), 
      .Q(\buffer[5][4][0] [15]), .QN());
   DFF_X1 \buffer_reg[5][4][0][14]  (.D(\input_filter[4][0] [14]), .CK(n_53_5), 
      .Q(\buffer[5][4][0] [14]), .QN());
   DFF_X1 \buffer_reg[5][4][0][13]  (.D(\input_filter[4][0] [13]), .CK(n_53_5), 
      .Q(\buffer[5][4][0] [13]), .QN());
   DFF_X1 \buffer_reg[5][4][0][12]  (.D(\input_filter[4][0] [12]), .CK(n_53_5), 
      .Q(\buffer[5][4][0] [12]), .QN());
   DFF_X1 \buffer_reg[5][4][0][11]  (.D(\input_filter[4][0] [11]), .CK(n_53_5), 
      .Q(\buffer[5][4][0] [11]), .QN());
   DFF_X1 \buffer_reg[5][4][0][10]  (.D(\input_filter[4][0] [10]), .CK(n_53_5), 
      .Q(\buffer[5][4][0] [10]), .QN());
   DFF_X1 \buffer_reg[5][4][0][9]  (.D(\input_filter[4][0] [9]), .CK(n_53_5), 
      .Q(\buffer[5][4][0] [9]), .QN());
   DFF_X1 \buffer_reg[5][4][0][8]  (.D(\input_filter[4][0] [8]), .CK(n_53_5), 
      .Q(\buffer[5][4][0] [8]), .QN());
   DFF_X1 \buffer_reg[5][4][0][7]  (.D(\input_filter[4][0] [7]), .CK(n_53_5), 
      .Q(\buffer[5][4][0] [7]), .QN());
   DFF_X1 \buffer_reg[5][4][0][6]  (.D(\input_filter[4][0] [6]), .CK(n_53_5), 
      .Q(\buffer[5][4][0] [6]), .QN());
   DFF_X1 \buffer_reg[5][4][0][5]  (.D(\input_filter[4][0] [5]), .CK(n_53_5), 
      .Q(\buffer[5][4][0] [5]), .QN());
   DFF_X1 \buffer_reg[5][4][0][4]  (.D(\input_filter[4][0] [4]), .CK(n_53_5), 
      .Q(\buffer[5][4][0] [4]), .QN());
   DFF_X1 \buffer_reg[5][4][0][3]  (.D(\input_filter[4][0] [3]), .CK(n_53_5), 
      .Q(\buffer[5][4][0] [3]), .QN());
   DFF_X1 \buffer_reg[5][4][0][2]  (.D(\input_filter[4][0] [2]), .CK(n_53_5), 
      .Q(\buffer[5][4][0] [2]), .QN());
   DFF_X1 \buffer_reg[5][4][0][1]  (.D(\input_filter[4][0] [1]), .CK(n_53_5), 
      .Q(\buffer[5][4][0] [1]), .QN());
   DFF_X1 \buffer_reg[5][4][0][0]  (.D(\input_filter[4][0] [0]), .CK(n_53_5), 
      .Q(\buffer[5][4][0] [0]), .QN());
   DFF_X1 \buffer_reg[4][4][0][15]  (.D(\input_filter[4][0] [15]), .CK(n_53_4), 
      .Q(\buffer[4][4][0] [15]), .QN());
   DFF_X1 \buffer_reg[4][4][0][14]  (.D(\input_filter[4][0] [14]), .CK(n_53_4), 
      .Q(\buffer[4][4][0] [14]), .QN());
   DFF_X1 \buffer_reg[4][4][0][13]  (.D(\input_filter[4][0] [13]), .CK(n_53_4), 
      .Q(\buffer[4][4][0] [13]), .QN());
   DFF_X1 \buffer_reg[4][4][0][12]  (.D(\input_filter[4][0] [12]), .CK(n_53_4), 
      .Q(\buffer[4][4][0] [12]), .QN());
   DFF_X1 \buffer_reg[4][4][0][11]  (.D(\input_filter[4][0] [11]), .CK(n_53_4), 
      .Q(\buffer[4][4][0] [11]), .QN());
   DFF_X1 \buffer_reg[4][4][0][10]  (.D(\input_filter[4][0] [10]), .CK(n_53_4), 
      .Q(\buffer[4][4][0] [10]), .QN());
   DFF_X1 \buffer_reg[4][4][0][9]  (.D(\input_filter[4][0] [9]), .CK(n_53_4), 
      .Q(\buffer[4][4][0] [9]), .QN());
   DFF_X1 \buffer_reg[4][4][0][8]  (.D(\input_filter[4][0] [8]), .CK(n_53_4), 
      .Q(\buffer[4][4][0] [8]), .QN());
   DFF_X1 \buffer_reg[4][4][0][7]  (.D(\input_filter[4][0] [7]), .CK(n_53_4), 
      .Q(\buffer[4][4][0] [7]), .QN());
   DFF_X1 \buffer_reg[4][4][0][6]  (.D(\input_filter[4][0] [6]), .CK(n_53_4), 
      .Q(\buffer[4][4][0] [6]), .QN());
   DFF_X1 \buffer_reg[4][4][0][5]  (.D(\input_filter[4][0] [5]), .CK(n_53_4), 
      .Q(\buffer[4][4][0] [5]), .QN());
   DFF_X1 \buffer_reg[4][4][0][4]  (.D(\input_filter[4][0] [4]), .CK(n_53_4), 
      .Q(\buffer[4][4][0] [4]), .QN());
   DFF_X1 \buffer_reg[4][4][0][3]  (.D(\input_filter[4][0] [3]), .CK(n_53_4), 
      .Q(\buffer[4][4][0] [3]), .QN());
   DFF_X1 \buffer_reg[4][4][0][2]  (.D(\input_filter[4][0] [2]), .CK(n_53_4), 
      .Q(\buffer[4][4][0] [2]), .QN());
   DFF_X1 \buffer_reg[4][4][0][1]  (.D(\input_filter[4][0] [1]), .CK(n_53_4), 
      .Q(\buffer[4][4][0] [1]), .QN());
   DFF_X1 \buffer_reg[4][4][0][0]  (.D(\input_filter[4][0] [0]), .CK(n_53_4), 
      .Q(\buffer[4][4][0] [0]), .QN());
   DFF_X1 \buffer_reg[3][4][0][15]  (.D(\input_filter[4][0] [15]), .CK(n_53_3), 
      .Q(\buffer[3][4][0] [15]), .QN());
   DFF_X1 \buffer_reg[3][4][0][14]  (.D(\input_filter[4][0] [14]), .CK(n_53_3), 
      .Q(\buffer[3][4][0] [14]), .QN());
   DFF_X1 \buffer_reg[3][4][0][13]  (.D(\input_filter[4][0] [13]), .CK(n_53_3), 
      .Q(\buffer[3][4][0] [13]), .QN());
   DFF_X1 \buffer_reg[3][4][0][12]  (.D(\input_filter[4][0] [12]), .CK(n_53_3), 
      .Q(\buffer[3][4][0] [12]), .QN());
   DFF_X1 \buffer_reg[3][4][0][11]  (.D(\input_filter[4][0] [11]), .CK(n_53_3), 
      .Q(\buffer[3][4][0] [11]), .QN());
   DFF_X1 \buffer_reg[3][4][0][10]  (.D(\input_filter[4][0] [10]), .CK(n_53_3), 
      .Q(\buffer[3][4][0] [10]), .QN());
   DFF_X1 \buffer_reg[3][4][0][9]  (.D(\input_filter[4][0] [9]), .CK(n_53_3), 
      .Q(\buffer[3][4][0] [9]), .QN());
   DFF_X1 \buffer_reg[3][4][0][8]  (.D(\input_filter[4][0] [8]), .CK(n_53_3), 
      .Q(\buffer[3][4][0] [8]), .QN());
   DFF_X1 \buffer_reg[3][4][0][7]  (.D(\input_filter[4][0] [7]), .CK(n_53_3), 
      .Q(\buffer[3][4][0] [7]), .QN());
   DFF_X1 \buffer_reg[3][4][0][6]  (.D(\input_filter[4][0] [6]), .CK(n_53_3), 
      .Q(\buffer[3][4][0] [6]), .QN());
   DFF_X1 \buffer_reg[3][4][0][5]  (.D(\input_filter[4][0] [5]), .CK(n_53_3), 
      .Q(\buffer[3][4][0] [5]), .QN());
   DFF_X1 \buffer_reg[3][4][0][4]  (.D(\input_filter[4][0] [4]), .CK(n_53_3), 
      .Q(\buffer[3][4][0] [4]), .QN());
   DFF_X1 \buffer_reg[3][4][0][3]  (.D(\input_filter[4][0] [3]), .CK(n_53_3), 
      .Q(\buffer[3][4][0] [3]), .QN());
   DFF_X1 \buffer_reg[3][4][0][2]  (.D(\input_filter[4][0] [2]), .CK(n_53_3), 
      .Q(\buffer[3][4][0] [2]), .QN());
   DFF_X1 \buffer_reg[3][4][0][1]  (.D(\input_filter[4][0] [1]), .CK(n_53_3), 
      .Q(\buffer[3][4][0] [1]), .QN());
   DFF_X1 \buffer_reg[3][4][0][0]  (.D(\input_filter[4][0] [0]), .CK(n_53_3), 
      .Q(\buffer[3][4][0] [0]), .QN());
   DFF_X1 \buffer_reg[2][4][0][15]  (.D(\input_filter[4][0] [15]), .CK(n_53_2), 
      .Q(\buffer[2][4][0] [15]), .QN());
   DFF_X1 \buffer_reg[2][4][0][14]  (.D(\input_filter[4][0] [14]), .CK(n_53_2), 
      .Q(\buffer[2][4][0] [14]), .QN());
   DFF_X1 \buffer_reg[2][4][0][13]  (.D(\input_filter[4][0] [13]), .CK(n_53_2), 
      .Q(\buffer[2][4][0] [13]), .QN());
   DFF_X1 \buffer_reg[2][4][0][12]  (.D(\input_filter[4][0] [12]), .CK(n_53_2), 
      .Q(\buffer[2][4][0] [12]), .QN());
   DFF_X1 \buffer_reg[2][4][0][11]  (.D(\input_filter[4][0] [11]), .CK(n_53_2), 
      .Q(\buffer[2][4][0] [11]), .QN());
   DFF_X1 \buffer_reg[2][4][0][10]  (.D(\input_filter[4][0] [10]), .CK(n_53_2), 
      .Q(\buffer[2][4][0] [10]), .QN());
   DFF_X1 \buffer_reg[2][4][0][9]  (.D(\input_filter[4][0] [9]), .CK(n_53_2), 
      .Q(\buffer[2][4][0] [9]), .QN());
   DFF_X1 \buffer_reg[2][4][0][8]  (.D(\input_filter[4][0] [8]), .CK(n_53_2), 
      .Q(\buffer[2][4][0] [8]), .QN());
   DFF_X1 \buffer_reg[2][4][0][7]  (.D(\input_filter[4][0] [7]), .CK(n_53_2), 
      .Q(\buffer[2][4][0] [7]), .QN());
   DFF_X1 \buffer_reg[2][4][0][6]  (.D(\input_filter[4][0] [6]), .CK(n_53_2), 
      .Q(\buffer[2][4][0] [6]), .QN());
   DFF_X1 \buffer_reg[2][4][0][5]  (.D(\input_filter[4][0] [5]), .CK(n_53_2), 
      .Q(\buffer[2][4][0] [5]), .QN());
   DFF_X1 \buffer_reg[2][4][0][4]  (.D(\input_filter[4][0] [4]), .CK(n_53_2), 
      .Q(\buffer[2][4][0] [4]), .QN());
   DFF_X1 \buffer_reg[2][4][0][3]  (.D(\input_filter[4][0] [3]), .CK(n_53_2), 
      .Q(\buffer[2][4][0] [3]), .QN());
   DFF_X1 \buffer_reg[2][4][0][2]  (.D(\input_filter[4][0] [2]), .CK(n_53_2), 
      .Q(\buffer[2][4][0] [2]), .QN());
   DFF_X1 \buffer_reg[2][4][0][1]  (.D(\input_filter[4][0] [1]), .CK(n_53_2), 
      .Q(\buffer[2][4][0] [1]), .QN());
   DFF_X1 \buffer_reg[2][4][0][0]  (.D(\input_filter[4][0] [0]), .CK(n_53_2), 
      .Q(\buffer[2][4][0] [0]), .QN());
   DFF_X1 \buffer_reg[1][4][0][15]  (.D(\input_filter[4][0] [15]), .CK(n_53_1), 
      .Q(\buffer[1][4][0] [15]), .QN());
   DFF_X1 \buffer_reg[1][4][0][14]  (.D(\input_filter[4][0] [14]), .CK(n_53_1), 
      .Q(\buffer[1][4][0] [14]), .QN());
   DFF_X1 \buffer_reg[1][4][0][13]  (.D(\input_filter[4][0] [13]), .CK(n_53_1), 
      .Q(\buffer[1][4][0] [13]), .QN());
   DFF_X1 \buffer_reg[1][4][0][12]  (.D(\input_filter[4][0] [12]), .CK(n_53_1), 
      .Q(\buffer[1][4][0] [12]), .QN());
   DFF_X1 \buffer_reg[1][4][0][11]  (.D(\input_filter[4][0] [11]), .CK(n_53_1), 
      .Q(\buffer[1][4][0] [11]), .QN());
   DFF_X1 \buffer_reg[1][4][0][10]  (.D(\input_filter[4][0] [10]), .CK(n_53_1), 
      .Q(\buffer[1][4][0] [10]), .QN());
   DFF_X1 \buffer_reg[1][4][0][9]  (.D(\input_filter[4][0] [9]), .CK(n_53_1), 
      .Q(\buffer[1][4][0] [9]), .QN());
   DFF_X1 \buffer_reg[1][4][0][8]  (.D(\input_filter[4][0] [8]), .CK(n_53_1), 
      .Q(\buffer[1][4][0] [8]), .QN());
   DFF_X1 \buffer_reg[1][4][0][7]  (.D(\input_filter[4][0] [7]), .CK(n_53_1), 
      .Q(\buffer[1][4][0] [7]), .QN());
   DFF_X1 \buffer_reg[1][4][0][6]  (.D(\input_filter[4][0] [6]), .CK(n_53_1), 
      .Q(\buffer[1][4][0] [6]), .QN());
   DFF_X1 \buffer_reg[1][4][0][5]  (.D(\input_filter[4][0] [5]), .CK(n_53_1), 
      .Q(\buffer[1][4][0] [5]), .QN());
   DFF_X1 \buffer_reg[1][4][0][4]  (.D(\input_filter[4][0] [4]), .CK(n_53_1), 
      .Q(\buffer[1][4][0] [4]), .QN());
   DFF_X1 \buffer_reg[1][4][0][3]  (.D(\input_filter[4][0] [3]), .CK(n_53_1), 
      .Q(\buffer[1][4][0] [3]), .QN());
   DFF_X1 \buffer_reg[1][4][0][2]  (.D(\input_filter[4][0] [2]), .CK(n_53_1), 
      .Q(\buffer[1][4][0] [2]), .QN());
   DFF_X1 \buffer_reg[1][4][0][1]  (.D(\input_filter[4][0] [1]), .CK(n_53_1), 
      .Q(\buffer[1][4][0] [1]), .QN());
   DFF_X1 \buffer_reg[1][4][0][0]  (.D(\input_filter[4][0] [0]), .CK(n_53_1), 
      .Q(\buffer[1][4][0] [0]), .QN());
   DFF_X1 \buffer_reg[0][4][0][15]  (.D(\input_filter[4][0] [15]), .CK(n_53_0), 
      .Q(\buffer[0][4][0] [15]), .QN());
   DFF_X1 \buffer_reg[0][4][0][14]  (.D(\input_filter[4][0] [14]), .CK(n_53_0), 
      .Q(\buffer[0][4][0] [14]), .QN());
   DFF_X1 \buffer_reg[0][4][0][13]  (.D(\input_filter[4][0] [13]), .CK(n_53_0), 
      .Q(\buffer[0][4][0] [13]), .QN());
   DFF_X1 \buffer_reg[0][4][0][12]  (.D(\input_filter[4][0] [12]), .CK(n_53_0), 
      .Q(\buffer[0][4][0] [12]), .QN());
   DFF_X1 \buffer_reg[0][4][0][11]  (.D(\input_filter[4][0] [11]), .CK(n_53_0), 
      .Q(\buffer[0][4][0] [11]), .QN());
   DFF_X1 \buffer_reg[0][4][0][10]  (.D(\input_filter[4][0] [10]), .CK(n_53_0), 
      .Q(\buffer[0][4][0] [10]), .QN());
   DFF_X1 \buffer_reg[0][4][0][9]  (.D(\input_filter[4][0] [9]), .CK(n_53_0), 
      .Q(\buffer[0][4][0] [9]), .QN());
   DFF_X1 \buffer_reg[0][4][0][8]  (.D(\input_filter[4][0] [8]), .CK(n_53_0), 
      .Q(\buffer[0][4][0] [8]), .QN());
   DFF_X1 \buffer_reg[0][4][0][7]  (.D(\input_filter[4][0] [7]), .CK(n_53_0), 
      .Q(\buffer[0][4][0] [7]), .QN());
   DFF_X1 \buffer_reg[0][4][0][6]  (.D(\input_filter[4][0] [6]), .CK(n_53_0), 
      .Q(\buffer[0][4][0] [6]), .QN());
   DFF_X1 \buffer_reg[0][4][0][5]  (.D(\input_filter[4][0] [5]), .CK(n_53_0), 
      .Q(\buffer[0][4][0] [5]), .QN());
   DFF_X1 \buffer_reg[0][4][0][4]  (.D(\input_filter[4][0] [4]), .CK(n_53_0), 
      .Q(\buffer[0][4][0] [4]), .QN());
   DFF_X1 \buffer_reg[0][4][0][3]  (.D(\input_filter[4][0] [3]), .CK(n_53_0), 
      .Q(\buffer[0][4][0] [3]), .QN());
   DFF_X1 \buffer_reg[0][4][0][2]  (.D(\input_filter[4][0] [2]), .CK(n_53_0), 
      .Q(\buffer[0][4][0] [2]), .QN());
   DFF_X1 \buffer_reg[0][4][0][1]  (.D(\input_filter[4][0] [1]), .CK(n_53_0), 
      .Q(\buffer[0][4][0] [1]), .QN());
   DFF_X1 \buffer_reg[0][4][0][0]  (.D(\input_filter[4][0] [0]), .CK(n_53_0), 
      .Q(\buffer[0][4][0] [0]), .QN());
   DFF_X1 \buffer_reg[15][3][4][15]  (.D(\input_filter[3][4] [15]), .CK(n_53_15), 
      .Q(\buffer[15][3][4] [15]), .QN());
   DFF_X1 \buffer_reg[15][3][4][14]  (.D(\input_filter[3][4] [14]), .CK(n_53_15), 
      .Q(\buffer[15][3][4] [14]), .QN());
   DFF_X1 \buffer_reg[15][3][4][13]  (.D(\input_filter[3][4] [13]), .CK(n_53_15), 
      .Q(\buffer[15][3][4] [13]), .QN());
   DFF_X1 \buffer_reg[15][3][4][12]  (.D(\input_filter[3][4] [12]), .CK(n_53_15), 
      .Q(\buffer[15][3][4] [12]), .QN());
   DFF_X1 \buffer_reg[15][3][4][11]  (.D(\input_filter[3][4] [11]), .CK(n_53_15), 
      .Q(\buffer[15][3][4] [11]), .QN());
   DFF_X1 \buffer_reg[15][3][4][10]  (.D(\input_filter[3][4] [10]), .CK(n_53_15), 
      .Q(\buffer[15][3][4] [10]), .QN());
   DFF_X1 \buffer_reg[15][3][4][9]  (.D(\input_filter[3][4] [9]), .CK(n_53_15), 
      .Q(\buffer[15][3][4] [9]), .QN());
   DFF_X1 \buffer_reg[15][3][4][8]  (.D(\input_filter[3][4] [8]), .CK(n_53_15), 
      .Q(\buffer[15][3][4] [8]), .QN());
   DFF_X1 \buffer_reg[15][3][4][7]  (.D(\input_filter[3][4] [7]), .CK(n_53_15), 
      .Q(\buffer[15][3][4] [7]), .QN());
   DFF_X1 \buffer_reg[15][3][4][6]  (.D(\input_filter[3][4] [6]), .CK(n_53_15), 
      .Q(\buffer[15][3][4] [6]), .QN());
   DFF_X1 \buffer_reg[15][3][4][5]  (.D(\input_filter[3][4] [5]), .CK(n_53_15), 
      .Q(\buffer[15][3][4] [5]), .QN());
   DFF_X1 \buffer_reg[15][3][4][4]  (.D(\input_filter[3][4] [4]), .CK(n_53_15), 
      .Q(\buffer[15][3][4] [4]), .QN());
   DFF_X1 \buffer_reg[15][3][4][3]  (.D(\input_filter[3][4] [3]), .CK(n_53_15), 
      .Q(\buffer[15][3][4] [3]), .QN());
   DFF_X1 \buffer_reg[15][3][4][2]  (.D(\input_filter[3][4] [2]), .CK(n_53_15), 
      .Q(\buffer[15][3][4] [2]), .QN());
   DFF_X1 \buffer_reg[15][3][4][1]  (.D(\input_filter[3][4] [1]), .CK(n_53_15), 
      .Q(\buffer[15][3][4] [1]), .QN());
   DFF_X1 \buffer_reg[15][3][4][0]  (.D(\input_filter[3][4] [0]), .CK(n_53_15), 
      .Q(\buffer[15][3][4] [0]), .QN());
   DFF_X1 \buffer_reg[14][3][4][15]  (.D(\input_filter[3][4] [15]), .CK(n_53_14), 
      .Q(\buffer[14][3][4] [15]), .QN());
   DFF_X1 \buffer_reg[14][3][4][14]  (.D(\input_filter[3][4] [14]), .CK(n_53_14), 
      .Q(\buffer[14][3][4] [14]), .QN());
   DFF_X1 \buffer_reg[14][3][4][13]  (.D(\input_filter[3][4] [13]), .CK(n_53_14), 
      .Q(\buffer[14][3][4] [13]), .QN());
   DFF_X1 \buffer_reg[14][3][4][12]  (.D(\input_filter[3][4] [12]), .CK(n_53_14), 
      .Q(\buffer[14][3][4] [12]), .QN());
   DFF_X1 \buffer_reg[14][3][4][11]  (.D(\input_filter[3][4] [11]), .CK(n_53_14), 
      .Q(\buffer[14][3][4] [11]), .QN());
   DFF_X1 \buffer_reg[14][3][4][10]  (.D(\input_filter[3][4] [10]), .CK(n_53_14), 
      .Q(\buffer[14][3][4] [10]), .QN());
   DFF_X1 \buffer_reg[14][3][4][9]  (.D(\input_filter[3][4] [9]), .CK(n_53_14), 
      .Q(\buffer[14][3][4] [9]), .QN());
   DFF_X1 \buffer_reg[14][3][4][8]  (.D(\input_filter[3][4] [8]), .CK(n_53_14), 
      .Q(\buffer[14][3][4] [8]), .QN());
   DFF_X1 \buffer_reg[14][3][4][7]  (.D(\input_filter[3][4] [7]), .CK(n_53_14), 
      .Q(\buffer[14][3][4] [7]), .QN());
   DFF_X1 \buffer_reg[14][3][4][6]  (.D(\input_filter[3][4] [6]), .CK(n_53_14), 
      .Q(\buffer[14][3][4] [6]), .QN());
   DFF_X1 \buffer_reg[14][3][4][5]  (.D(\input_filter[3][4] [5]), .CK(n_53_14), 
      .Q(\buffer[14][3][4] [5]), .QN());
   DFF_X1 \buffer_reg[14][3][4][4]  (.D(\input_filter[3][4] [4]), .CK(n_53_14), 
      .Q(\buffer[14][3][4] [4]), .QN());
   DFF_X1 \buffer_reg[14][3][4][3]  (.D(\input_filter[3][4] [3]), .CK(n_53_14), 
      .Q(\buffer[14][3][4] [3]), .QN());
   DFF_X1 \buffer_reg[14][3][4][2]  (.D(\input_filter[3][4] [2]), .CK(n_53_14), 
      .Q(\buffer[14][3][4] [2]), .QN());
   DFF_X1 \buffer_reg[14][3][4][1]  (.D(\input_filter[3][4] [1]), .CK(n_53_14), 
      .Q(\buffer[14][3][4] [1]), .QN());
   DFF_X1 \buffer_reg[14][3][4][0]  (.D(\input_filter[3][4] [0]), .CK(n_53_14), 
      .Q(\buffer[14][3][4] [0]), .QN());
   DFF_X1 \buffer_reg[13][3][4][15]  (.D(\input_filter[3][4] [15]), .CK(n_53_13), 
      .Q(\buffer[13][3][4] [15]), .QN());
   DFF_X1 \buffer_reg[13][3][4][14]  (.D(\input_filter[3][4] [14]), .CK(n_53_13), 
      .Q(\buffer[13][3][4] [14]), .QN());
   DFF_X1 \buffer_reg[13][3][4][13]  (.D(\input_filter[3][4] [13]), .CK(n_53_13), 
      .Q(\buffer[13][3][4] [13]), .QN());
   DFF_X1 \buffer_reg[13][3][4][12]  (.D(\input_filter[3][4] [12]), .CK(n_53_13), 
      .Q(\buffer[13][3][4] [12]), .QN());
   DFF_X1 \buffer_reg[13][3][4][11]  (.D(\input_filter[3][4] [11]), .CK(n_53_13), 
      .Q(\buffer[13][3][4] [11]), .QN());
   DFF_X1 \buffer_reg[13][3][4][10]  (.D(\input_filter[3][4] [10]), .CK(n_53_13), 
      .Q(\buffer[13][3][4] [10]), .QN());
   DFF_X1 \buffer_reg[13][3][4][9]  (.D(\input_filter[3][4] [9]), .CK(n_53_13), 
      .Q(\buffer[13][3][4] [9]), .QN());
   DFF_X1 \buffer_reg[13][3][4][8]  (.D(\input_filter[3][4] [8]), .CK(n_53_13), 
      .Q(\buffer[13][3][4] [8]), .QN());
   DFF_X1 \buffer_reg[13][3][4][7]  (.D(\input_filter[3][4] [7]), .CK(n_53_13), 
      .Q(\buffer[13][3][4] [7]), .QN());
   DFF_X1 \buffer_reg[13][3][4][6]  (.D(\input_filter[3][4] [6]), .CK(n_53_13), 
      .Q(\buffer[13][3][4] [6]), .QN());
   DFF_X1 \buffer_reg[13][3][4][5]  (.D(\input_filter[3][4] [5]), .CK(n_53_13), 
      .Q(\buffer[13][3][4] [5]), .QN());
   DFF_X1 \buffer_reg[13][3][4][4]  (.D(\input_filter[3][4] [4]), .CK(n_53_13), 
      .Q(\buffer[13][3][4] [4]), .QN());
   DFF_X1 \buffer_reg[13][3][4][3]  (.D(\input_filter[3][4] [3]), .CK(n_53_13), 
      .Q(\buffer[13][3][4] [3]), .QN());
   DFF_X1 \buffer_reg[13][3][4][2]  (.D(\input_filter[3][4] [2]), .CK(n_53_13), 
      .Q(\buffer[13][3][4] [2]), .QN());
   DFF_X1 \buffer_reg[13][3][4][1]  (.D(\input_filter[3][4] [1]), .CK(n_53_13), 
      .Q(\buffer[13][3][4] [1]), .QN());
   DFF_X1 \buffer_reg[13][3][4][0]  (.D(\input_filter[3][4] [0]), .CK(n_53_13), 
      .Q(\buffer[13][3][4] [0]), .QN());
   DFF_X1 \buffer_reg[12][3][4][15]  (.D(\input_filter[3][4] [15]), .CK(n_53_12), 
      .Q(\buffer[12][3][4] [15]), .QN());
   DFF_X1 \buffer_reg[12][3][4][14]  (.D(\input_filter[3][4] [14]), .CK(n_53_12), 
      .Q(\buffer[12][3][4] [14]), .QN());
   DFF_X1 \buffer_reg[12][3][4][13]  (.D(\input_filter[3][4] [13]), .CK(n_53_12), 
      .Q(\buffer[12][3][4] [13]), .QN());
   DFF_X1 \buffer_reg[12][3][4][12]  (.D(\input_filter[3][4] [12]), .CK(n_53_12), 
      .Q(\buffer[12][3][4] [12]), .QN());
   DFF_X1 \buffer_reg[12][3][4][11]  (.D(\input_filter[3][4] [11]), .CK(n_53_12), 
      .Q(\buffer[12][3][4] [11]), .QN());
   DFF_X1 \buffer_reg[12][3][4][10]  (.D(\input_filter[3][4] [10]), .CK(n_53_12), 
      .Q(\buffer[12][3][4] [10]), .QN());
   DFF_X1 \buffer_reg[12][3][4][9]  (.D(\input_filter[3][4] [9]), .CK(n_53_12), 
      .Q(\buffer[12][3][4] [9]), .QN());
   DFF_X1 \buffer_reg[12][3][4][8]  (.D(\input_filter[3][4] [8]), .CK(n_53_12), 
      .Q(\buffer[12][3][4] [8]), .QN());
   DFF_X1 \buffer_reg[12][3][4][7]  (.D(\input_filter[3][4] [7]), .CK(n_53_12), 
      .Q(\buffer[12][3][4] [7]), .QN());
   DFF_X1 \buffer_reg[12][3][4][6]  (.D(\input_filter[3][4] [6]), .CK(n_53_12), 
      .Q(\buffer[12][3][4] [6]), .QN());
   DFF_X1 \buffer_reg[12][3][4][5]  (.D(\input_filter[3][4] [5]), .CK(n_53_12), 
      .Q(\buffer[12][3][4] [5]), .QN());
   DFF_X1 \buffer_reg[12][3][4][4]  (.D(\input_filter[3][4] [4]), .CK(n_53_12), 
      .Q(\buffer[12][3][4] [4]), .QN());
   DFF_X1 \buffer_reg[12][3][4][3]  (.D(\input_filter[3][4] [3]), .CK(n_53_12), 
      .Q(\buffer[12][3][4] [3]), .QN());
   DFF_X1 \buffer_reg[12][3][4][2]  (.D(\input_filter[3][4] [2]), .CK(n_53_12), 
      .Q(\buffer[12][3][4] [2]), .QN());
   DFF_X1 \buffer_reg[12][3][4][1]  (.D(\input_filter[3][4] [1]), .CK(n_53_12), 
      .Q(\buffer[12][3][4] [1]), .QN());
   DFF_X1 \buffer_reg[12][3][4][0]  (.D(\input_filter[3][4] [0]), .CK(n_53_12), 
      .Q(\buffer[12][3][4] [0]), .QN());
   DFF_X1 \buffer_reg[11][3][4][15]  (.D(\input_filter[3][4] [15]), .CK(n_53_11), 
      .Q(\buffer[11][3][4] [15]), .QN());
   DFF_X1 \buffer_reg[11][3][4][14]  (.D(\input_filter[3][4] [14]), .CK(n_53_11), 
      .Q(\buffer[11][3][4] [14]), .QN());
   DFF_X1 \buffer_reg[11][3][4][13]  (.D(\input_filter[3][4] [13]), .CK(n_53_11), 
      .Q(\buffer[11][3][4] [13]), .QN());
   DFF_X1 \buffer_reg[11][3][4][12]  (.D(\input_filter[3][4] [12]), .CK(n_53_11), 
      .Q(\buffer[11][3][4] [12]), .QN());
   DFF_X1 \buffer_reg[11][3][4][11]  (.D(\input_filter[3][4] [11]), .CK(n_53_11), 
      .Q(\buffer[11][3][4] [11]), .QN());
   DFF_X1 \buffer_reg[11][3][4][10]  (.D(\input_filter[3][4] [10]), .CK(n_53_11), 
      .Q(\buffer[11][3][4] [10]), .QN());
   DFF_X1 \buffer_reg[11][3][4][9]  (.D(\input_filter[3][4] [9]), .CK(n_53_11), 
      .Q(\buffer[11][3][4] [9]), .QN());
   DFF_X1 \buffer_reg[11][3][4][8]  (.D(\input_filter[3][4] [8]), .CK(n_53_11), 
      .Q(\buffer[11][3][4] [8]), .QN());
   DFF_X1 \buffer_reg[11][3][4][7]  (.D(\input_filter[3][4] [7]), .CK(n_53_11), 
      .Q(\buffer[11][3][4] [7]), .QN());
   DFF_X1 \buffer_reg[11][3][4][6]  (.D(\input_filter[3][4] [6]), .CK(n_53_11), 
      .Q(\buffer[11][3][4] [6]), .QN());
   DFF_X1 \buffer_reg[11][3][4][5]  (.D(\input_filter[3][4] [5]), .CK(n_53_11), 
      .Q(\buffer[11][3][4] [5]), .QN());
   DFF_X1 \buffer_reg[11][3][4][4]  (.D(\input_filter[3][4] [4]), .CK(n_53_11), 
      .Q(\buffer[11][3][4] [4]), .QN());
   DFF_X1 \buffer_reg[11][3][4][3]  (.D(\input_filter[3][4] [3]), .CK(n_53_11), 
      .Q(\buffer[11][3][4] [3]), .QN());
   DFF_X1 \buffer_reg[11][3][4][2]  (.D(\input_filter[3][4] [2]), .CK(n_53_11), 
      .Q(\buffer[11][3][4] [2]), .QN());
   DFF_X1 \buffer_reg[11][3][4][1]  (.D(\input_filter[3][4] [1]), .CK(n_53_11), 
      .Q(\buffer[11][3][4] [1]), .QN());
   DFF_X1 \buffer_reg[11][3][4][0]  (.D(\input_filter[3][4] [0]), .CK(n_53_11), 
      .Q(\buffer[11][3][4] [0]), .QN());
   DFF_X1 \buffer_reg[10][3][4][15]  (.D(\input_filter[3][4] [15]), .CK(n_53_10), 
      .Q(\buffer[10][3][4] [15]), .QN());
   DFF_X1 \buffer_reg[10][3][4][14]  (.D(\input_filter[3][4] [14]), .CK(n_53_10), 
      .Q(\buffer[10][3][4] [14]), .QN());
   DFF_X1 \buffer_reg[10][3][4][13]  (.D(\input_filter[3][4] [13]), .CK(n_53_10), 
      .Q(\buffer[10][3][4] [13]), .QN());
   DFF_X1 \buffer_reg[10][3][4][12]  (.D(\input_filter[3][4] [12]), .CK(n_53_10), 
      .Q(\buffer[10][3][4] [12]), .QN());
   DFF_X1 \buffer_reg[10][3][4][11]  (.D(\input_filter[3][4] [11]), .CK(n_53_10), 
      .Q(\buffer[10][3][4] [11]), .QN());
   DFF_X1 \buffer_reg[10][3][4][10]  (.D(\input_filter[3][4] [10]), .CK(n_53_10), 
      .Q(\buffer[10][3][4] [10]), .QN());
   DFF_X1 \buffer_reg[10][3][4][9]  (.D(\input_filter[3][4] [9]), .CK(n_53_10), 
      .Q(\buffer[10][3][4] [9]), .QN());
   DFF_X1 \buffer_reg[10][3][4][8]  (.D(\input_filter[3][4] [8]), .CK(n_53_10), 
      .Q(\buffer[10][3][4] [8]), .QN());
   DFF_X1 \buffer_reg[10][3][4][7]  (.D(\input_filter[3][4] [7]), .CK(n_53_10), 
      .Q(\buffer[10][3][4] [7]), .QN());
   DFF_X1 \buffer_reg[10][3][4][6]  (.D(\input_filter[3][4] [6]), .CK(n_53_10), 
      .Q(\buffer[10][3][4] [6]), .QN());
   DFF_X1 \buffer_reg[10][3][4][5]  (.D(\input_filter[3][4] [5]), .CK(n_53_10), 
      .Q(\buffer[10][3][4] [5]), .QN());
   DFF_X1 \buffer_reg[10][3][4][4]  (.D(\input_filter[3][4] [4]), .CK(n_53_10), 
      .Q(\buffer[10][3][4] [4]), .QN());
   DFF_X1 \buffer_reg[10][3][4][3]  (.D(\input_filter[3][4] [3]), .CK(n_53_10), 
      .Q(\buffer[10][3][4] [3]), .QN());
   DFF_X1 \buffer_reg[10][3][4][2]  (.D(\input_filter[3][4] [2]), .CK(n_53_10), 
      .Q(\buffer[10][3][4] [2]), .QN());
   DFF_X1 \buffer_reg[10][3][4][1]  (.D(\input_filter[3][4] [1]), .CK(n_53_10), 
      .Q(\buffer[10][3][4] [1]), .QN());
   DFF_X1 \buffer_reg[10][3][4][0]  (.D(\input_filter[3][4] [0]), .CK(n_53_10), 
      .Q(\buffer[10][3][4] [0]), .QN());
   DFF_X1 \buffer_reg[9][3][4][15]  (.D(\input_filter[3][4] [15]), .CK(n_53_9), 
      .Q(\buffer[9][3][4] [15]), .QN());
   DFF_X1 \buffer_reg[9][3][4][14]  (.D(\input_filter[3][4] [14]), .CK(n_53_9), 
      .Q(\buffer[9][3][4] [14]), .QN());
   DFF_X1 \buffer_reg[9][3][4][13]  (.D(\input_filter[3][4] [13]), .CK(n_53_9), 
      .Q(\buffer[9][3][4] [13]), .QN());
   DFF_X1 \buffer_reg[9][3][4][12]  (.D(\input_filter[3][4] [12]), .CK(n_53_9), 
      .Q(\buffer[9][3][4] [12]), .QN());
   DFF_X1 \buffer_reg[9][3][4][11]  (.D(\input_filter[3][4] [11]), .CK(n_53_9), 
      .Q(\buffer[9][3][4] [11]), .QN());
   DFF_X1 \buffer_reg[9][3][4][10]  (.D(\input_filter[3][4] [10]), .CK(n_53_9), 
      .Q(\buffer[9][3][4] [10]), .QN());
   DFF_X1 \buffer_reg[9][3][4][9]  (.D(\input_filter[3][4] [9]), .CK(n_53_9), 
      .Q(\buffer[9][3][4] [9]), .QN());
   DFF_X1 \buffer_reg[9][3][4][8]  (.D(\input_filter[3][4] [8]), .CK(n_53_9), 
      .Q(\buffer[9][3][4] [8]), .QN());
   DFF_X1 \buffer_reg[9][3][4][7]  (.D(\input_filter[3][4] [7]), .CK(n_53_9), 
      .Q(\buffer[9][3][4] [7]), .QN());
   DFF_X1 \buffer_reg[9][3][4][6]  (.D(\input_filter[3][4] [6]), .CK(n_53_9), 
      .Q(\buffer[9][3][4] [6]), .QN());
   DFF_X1 \buffer_reg[9][3][4][5]  (.D(\input_filter[3][4] [5]), .CK(n_53_9), 
      .Q(\buffer[9][3][4] [5]), .QN());
   DFF_X1 \buffer_reg[9][3][4][4]  (.D(\input_filter[3][4] [4]), .CK(n_53_9), 
      .Q(\buffer[9][3][4] [4]), .QN());
   DFF_X1 \buffer_reg[9][3][4][3]  (.D(\input_filter[3][4] [3]), .CK(n_53_9), 
      .Q(\buffer[9][3][4] [3]), .QN());
   DFF_X1 \buffer_reg[9][3][4][2]  (.D(\input_filter[3][4] [2]), .CK(n_53_9), 
      .Q(\buffer[9][3][4] [2]), .QN());
   DFF_X1 \buffer_reg[9][3][4][1]  (.D(\input_filter[3][4] [1]), .CK(n_53_9), 
      .Q(\buffer[9][3][4] [1]), .QN());
   DFF_X1 \buffer_reg[9][3][4][0]  (.D(\input_filter[3][4] [0]), .CK(n_53_9), 
      .Q(\buffer[9][3][4] [0]), .QN());
   DFF_X1 \buffer_reg[8][3][4][15]  (.D(\input_filter[3][4] [15]), .CK(n_53_8), 
      .Q(\buffer[8][3][4] [15]), .QN());
   DFF_X1 \buffer_reg[8][3][4][14]  (.D(\input_filter[3][4] [14]), .CK(n_53_8), 
      .Q(\buffer[8][3][4] [14]), .QN());
   DFF_X1 \buffer_reg[8][3][4][13]  (.D(\input_filter[3][4] [13]), .CK(n_53_8), 
      .Q(\buffer[8][3][4] [13]), .QN());
   DFF_X1 \buffer_reg[8][3][4][12]  (.D(\input_filter[3][4] [12]), .CK(n_53_8), 
      .Q(\buffer[8][3][4] [12]), .QN());
   DFF_X1 \buffer_reg[8][3][4][11]  (.D(\input_filter[3][4] [11]), .CK(n_53_8), 
      .Q(\buffer[8][3][4] [11]), .QN());
   DFF_X1 \buffer_reg[8][3][4][10]  (.D(\input_filter[3][4] [10]), .CK(n_53_8), 
      .Q(\buffer[8][3][4] [10]), .QN());
   DFF_X1 \buffer_reg[8][3][4][9]  (.D(\input_filter[3][4] [9]), .CK(n_53_8), 
      .Q(\buffer[8][3][4] [9]), .QN());
   DFF_X1 \buffer_reg[8][3][4][8]  (.D(\input_filter[3][4] [8]), .CK(n_53_8), 
      .Q(\buffer[8][3][4] [8]), .QN());
   DFF_X1 \buffer_reg[8][3][4][7]  (.D(\input_filter[3][4] [7]), .CK(n_53_8), 
      .Q(\buffer[8][3][4] [7]), .QN());
   DFF_X1 \buffer_reg[8][3][4][6]  (.D(\input_filter[3][4] [6]), .CK(n_53_8), 
      .Q(\buffer[8][3][4] [6]), .QN());
   DFF_X1 \buffer_reg[8][3][4][5]  (.D(\input_filter[3][4] [5]), .CK(n_53_8), 
      .Q(\buffer[8][3][4] [5]), .QN());
   DFF_X1 \buffer_reg[8][3][4][4]  (.D(\input_filter[3][4] [4]), .CK(n_53_8), 
      .Q(\buffer[8][3][4] [4]), .QN());
   DFF_X1 \buffer_reg[8][3][4][3]  (.D(\input_filter[3][4] [3]), .CK(n_53_8), 
      .Q(\buffer[8][3][4] [3]), .QN());
   DFF_X1 \buffer_reg[8][3][4][2]  (.D(\input_filter[3][4] [2]), .CK(n_53_8), 
      .Q(\buffer[8][3][4] [2]), .QN());
   DFF_X1 \buffer_reg[8][3][4][1]  (.D(\input_filter[3][4] [1]), .CK(n_53_8), 
      .Q(\buffer[8][3][4] [1]), .QN());
   DFF_X1 \buffer_reg[8][3][4][0]  (.D(\input_filter[3][4] [0]), .CK(n_53_8), 
      .Q(\buffer[8][3][4] [0]), .QN());
   DFF_X1 \buffer_reg[7][3][4][15]  (.D(\input_filter[3][4] [15]), .CK(n_53_7), 
      .Q(\buffer[7][3][4] [15]), .QN());
   DFF_X1 \buffer_reg[7][3][4][14]  (.D(\input_filter[3][4] [14]), .CK(n_53_7), 
      .Q(\buffer[7][3][4] [14]), .QN());
   DFF_X1 \buffer_reg[7][3][4][13]  (.D(\input_filter[3][4] [13]), .CK(n_53_7), 
      .Q(\buffer[7][3][4] [13]), .QN());
   DFF_X1 \buffer_reg[7][3][4][12]  (.D(\input_filter[3][4] [12]), .CK(n_53_7), 
      .Q(\buffer[7][3][4] [12]), .QN());
   DFF_X1 \buffer_reg[7][3][4][11]  (.D(\input_filter[3][4] [11]), .CK(n_53_7), 
      .Q(\buffer[7][3][4] [11]), .QN());
   DFF_X1 \buffer_reg[7][3][4][10]  (.D(\input_filter[3][4] [10]), .CK(n_53_7), 
      .Q(\buffer[7][3][4] [10]), .QN());
   DFF_X1 \buffer_reg[7][3][4][9]  (.D(\input_filter[3][4] [9]), .CK(n_53_7), 
      .Q(\buffer[7][3][4] [9]), .QN());
   DFF_X1 \buffer_reg[7][3][4][8]  (.D(\input_filter[3][4] [8]), .CK(n_53_7), 
      .Q(\buffer[7][3][4] [8]), .QN());
   DFF_X1 \buffer_reg[7][3][4][7]  (.D(\input_filter[3][4] [7]), .CK(n_53_7), 
      .Q(\buffer[7][3][4] [7]), .QN());
   DFF_X1 \buffer_reg[7][3][4][6]  (.D(\input_filter[3][4] [6]), .CK(n_53_7), 
      .Q(\buffer[7][3][4] [6]), .QN());
   DFF_X1 \buffer_reg[7][3][4][5]  (.D(\input_filter[3][4] [5]), .CK(n_53_7), 
      .Q(\buffer[7][3][4] [5]), .QN());
   DFF_X1 \buffer_reg[7][3][4][4]  (.D(\input_filter[3][4] [4]), .CK(n_53_7), 
      .Q(\buffer[7][3][4] [4]), .QN());
   DFF_X1 \buffer_reg[7][3][4][3]  (.D(\input_filter[3][4] [3]), .CK(n_53_7), 
      .Q(\buffer[7][3][4] [3]), .QN());
   DFF_X1 \buffer_reg[7][3][4][2]  (.D(\input_filter[3][4] [2]), .CK(n_53_7), 
      .Q(\buffer[7][3][4] [2]), .QN());
   DFF_X1 \buffer_reg[7][3][4][1]  (.D(\input_filter[3][4] [1]), .CK(n_53_7), 
      .Q(\buffer[7][3][4] [1]), .QN());
   DFF_X1 \buffer_reg[7][3][4][0]  (.D(\input_filter[3][4] [0]), .CK(n_53_7), 
      .Q(\buffer[7][3][4] [0]), .QN());
   DFF_X1 \buffer_reg[6][3][4][15]  (.D(\input_filter[3][4] [15]), .CK(n_53_6), 
      .Q(\buffer[6][3][4] [15]), .QN());
   DFF_X1 \buffer_reg[6][3][4][14]  (.D(\input_filter[3][4] [14]), .CK(n_53_6), 
      .Q(\buffer[6][3][4] [14]), .QN());
   DFF_X1 \buffer_reg[6][3][4][13]  (.D(\input_filter[3][4] [13]), .CK(n_53_6), 
      .Q(\buffer[6][3][4] [13]), .QN());
   DFF_X1 \buffer_reg[6][3][4][12]  (.D(\input_filter[3][4] [12]), .CK(n_53_6), 
      .Q(\buffer[6][3][4] [12]), .QN());
   DFF_X1 \buffer_reg[6][3][4][11]  (.D(\input_filter[3][4] [11]), .CK(n_53_6), 
      .Q(\buffer[6][3][4] [11]), .QN());
   DFF_X1 \buffer_reg[6][3][4][10]  (.D(\input_filter[3][4] [10]), .CK(n_53_6), 
      .Q(\buffer[6][3][4] [10]), .QN());
   DFF_X1 \buffer_reg[6][3][4][9]  (.D(\input_filter[3][4] [9]), .CK(n_53_6), 
      .Q(\buffer[6][3][4] [9]), .QN());
   DFF_X1 \buffer_reg[6][3][4][8]  (.D(\input_filter[3][4] [8]), .CK(n_53_6), 
      .Q(\buffer[6][3][4] [8]), .QN());
   DFF_X1 \buffer_reg[6][3][4][7]  (.D(\input_filter[3][4] [7]), .CK(n_53_6), 
      .Q(\buffer[6][3][4] [7]), .QN());
   DFF_X1 \buffer_reg[6][3][4][6]  (.D(\input_filter[3][4] [6]), .CK(n_53_6), 
      .Q(\buffer[6][3][4] [6]), .QN());
   DFF_X1 \buffer_reg[6][3][4][5]  (.D(\input_filter[3][4] [5]), .CK(n_53_6), 
      .Q(\buffer[6][3][4] [5]), .QN());
   DFF_X1 \buffer_reg[6][3][4][4]  (.D(\input_filter[3][4] [4]), .CK(n_53_6), 
      .Q(\buffer[6][3][4] [4]), .QN());
   DFF_X1 \buffer_reg[6][3][4][3]  (.D(\input_filter[3][4] [3]), .CK(n_53_6), 
      .Q(\buffer[6][3][4] [3]), .QN());
   DFF_X1 \buffer_reg[6][3][4][2]  (.D(\input_filter[3][4] [2]), .CK(n_53_6), 
      .Q(\buffer[6][3][4] [2]), .QN());
   DFF_X1 \buffer_reg[6][3][4][1]  (.D(\input_filter[3][4] [1]), .CK(n_53_6), 
      .Q(\buffer[6][3][4] [1]), .QN());
   DFF_X1 \buffer_reg[6][3][4][0]  (.D(\input_filter[3][4] [0]), .CK(n_53_6), 
      .Q(\buffer[6][3][4] [0]), .QN());
   CLKGATETST_X1 \clk_gate_buffer_reg[0][3][3]_reg  (.CK(read), .E(n_0), 
      .SE(1'b0), .GCK(n_53_0));
   CLKGATETST_X1 \clk_gate_buffer_reg[1][3][3]_reg  (.CK(read), .E(n_1), 
      .SE(1'b0), .GCK(n_53_1));
   CLKGATETST_X1 \clk_gate_buffer_reg[2][3][3]_reg  (.CK(read), .E(n_2), 
      .SE(1'b0), .GCK(n_53_2));
   CLKGATETST_X1 \clk_gate_buffer_reg[3][3][3]_reg  (.CK(read), .E(n_3), 
      .SE(1'b0), .GCK(n_53_3));
   CLKGATETST_X1 \clk_gate_buffer_reg[4][3][3]_reg  (.CK(read), .E(n_4), 
      .SE(1'b0), .GCK(n_53_4));
   CLKGATETST_X1 \clk_gate_buffer_reg[5][3][3]_reg  (.CK(read), .E(n_5), 
      .SE(1'b0), .GCK(n_53_5));
   CLKGATETST_X1 \clk_gate_buffer_reg[6][3][3]_reg  (.CK(read), .E(n_6), 
      .SE(1'b0), .GCK(n_53_6));
   CLKGATETST_X1 \clk_gate_buffer_reg[7][3][3]_reg  (.CK(read), .E(n_7), 
      .SE(1'b0), .GCK(n_53_7));
   CLKGATETST_X1 \clk_gate_buffer_reg[8][3][3]_reg  (.CK(read), .E(n_8), 
      .SE(1'b0), .GCK(n_53_8));
   CLKGATETST_X1 \clk_gate_buffer_reg[9][3][3]_reg  (.CK(read), .E(n_9), 
      .SE(1'b0), .GCK(n_53_9));
   CLKGATETST_X1 \clk_gate_buffer_reg[10][3][3]_reg  (.CK(read), .E(n_10), 
      .SE(1'b0), .GCK(n_53_10));
   CLKGATETST_X1 \clk_gate_buffer_reg[11][3][3]_reg  (.CK(read), .E(n_11), 
      .SE(1'b0), .GCK(n_53_11));
   CLKGATETST_X1 \clk_gate_buffer_reg[12][3][3]_reg  (.CK(read), .E(n_12), 
      .SE(1'b0), .GCK(n_53_12));
   CLKGATETST_X1 \clk_gate_buffer_reg[13][3][3]_reg  (.CK(read), .E(n_13), 
      .SE(1'b0), .GCK(n_53_13));
   CLKGATETST_X1 \clk_gate_buffer_reg[14][3][3]_reg  (.CK(read), .E(n_14), 
      .SE(1'b0), .GCK(n_53_14));
   CLKGATETST_X1 \clk_gate_buffer_reg[15][3][3]_reg  (.CK(read), .E(n_15), 
      .SE(1'b0), .GCK(n_53_15));
   DFF_X1 \buffer_reg[1][4][3][15]  (.D(\input_filter[4][3] [15]), .CK(n_54_3), 
      .Q(\buffer[1][4][3] [15]), .QN());
   DFF_X1 \buffer_reg[1][4][3][14]  (.D(\input_filter[4][3] [14]), .CK(n_54_3), 
      .Q(\buffer[1][4][3] [14]), .QN());
   DFF_X1 \buffer_reg[1][4][3][13]  (.D(\input_filter[4][3] [13]), .CK(n_54_3), 
      .Q(\buffer[1][4][3] [13]), .QN());
   DFF_X1 \buffer_reg[1][4][3][12]  (.D(\input_filter[4][3] [12]), .CK(n_54_3), 
      .Q(\buffer[1][4][3] [12]), .QN());
   DFF_X1 \buffer_reg[1][4][3][11]  (.D(\input_filter[4][3] [11]), .CK(n_54_3), 
      .Q(\buffer[1][4][3] [11]), .QN());
   DFF_X1 \buffer_reg[1][4][3][10]  (.D(\input_filter[4][3] [10]), .CK(n_54_3), 
      .Q(\buffer[1][4][3] [10]), .QN());
   DFF_X1 \buffer_reg[1][4][3][9]  (.D(\input_filter[4][3] [9]), .CK(n_54_3), 
      .Q(\buffer[1][4][3] [9]), .QN());
   DFF_X1 \buffer_reg[1][4][3][8]  (.D(\input_filter[4][3] [8]), .CK(n_54_3), 
      .Q(\buffer[1][4][3] [8]), .QN());
   DFF_X1 \buffer_reg[1][4][3][7]  (.D(\input_filter[4][3] [7]), .CK(n_54_3), 
      .Q(\buffer[1][4][3] [7]), .QN());
   DFF_X1 \buffer_reg[1][4][3][6]  (.D(\input_filter[4][3] [6]), .CK(n_54_3), 
      .Q(\buffer[1][4][3] [6]), .QN());
   DFF_X1 \buffer_reg[1][4][3][5]  (.D(\input_filter[4][3] [5]), .CK(n_54_3), 
      .Q(\buffer[1][4][3] [5]), .QN());
   DFF_X1 \buffer_reg[1][4][3][4]  (.D(\input_filter[4][3] [4]), .CK(n_54_3), 
      .Q(\buffer[1][4][3] [4]), .QN());
   DFF_X1 \buffer_reg[1][4][3][3]  (.D(\input_filter[4][3] [3]), .CK(n_54_3), 
      .Q(\buffer[1][4][3] [3]), .QN());
   DFF_X1 \buffer_reg[1][4][3][2]  (.D(\input_filter[4][3] [2]), .CK(n_54_3), 
      .Q(\buffer[1][4][3] [2]), .QN());
   DFF_X1 \buffer_reg[1][4][3][1]  (.D(\input_filter[4][3] [1]), .CK(n_54_3), 
      .Q(\buffer[1][4][3] [1]), .QN());
   DFF_X1 \buffer_reg[1][4][3][0]  (.D(\input_filter[4][3] [0]), .CK(n_54_3), 
      .Q(\buffer[1][4][3] [0]), .QN());
   DFF_X1 \buffer_reg[2][4][3][15]  (.D(\input_filter[4][3] [15]), .CK(n_54_4), 
      .Q(\buffer[2][4][3] [15]), .QN());
   DFF_X1 \buffer_reg[2][4][3][14]  (.D(\input_filter[4][3] [14]), .CK(n_54_4), 
      .Q(\buffer[2][4][3] [14]), .QN());
   DFF_X1 \buffer_reg[2][4][3][13]  (.D(\input_filter[4][3] [13]), .CK(n_54_4), 
      .Q(\buffer[2][4][3] [13]), .QN());
   DFF_X1 \buffer_reg[2][4][3][12]  (.D(\input_filter[4][3] [12]), .CK(n_54_4), 
      .Q(\buffer[2][4][3] [12]), .QN());
   DFF_X1 \buffer_reg[2][4][3][11]  (.D(\input_filter[4][3] [11]), .CK(n_54_4), 
      .Q(\buffer[2][4][3] [11]), .QN());
   DFF_X1 \buffer_reg[2][4][3][10]  (.D(\input_filter[4][3] [10]), .CK(n_54_4), 
      .Q(\buffer[2][4][3] [10]), .QN());
   DFF_X1 \buffer_reg[2][4][3][9]  (.D(\input_filter[4][3] [9]), .CK(n_54_4), 
      .Q(\buffer[2][4][3] [9]), .QN());
   DFF_X1 \buffer_reg[2][4][3][8]  (.D(\input_filter[4][3] [8]), .CK(n_54_4), 
      .Q(\buffer[2][4][3] [8]), .QN());
   DFF_X1 \buffer_reg[2][4][3][7]  (.D(\input_filter[4][3] [7]), .CK(n_54_4), 
      .Q(\buffer[2][4][3] [7]), .QN());
   DFF_X1 \buffer_reg[2][4][3][6]  (.D(\input_filter[4][3] [6]), .CK(n_54_4), 
      .Q(\buffer[2][4][3] [6]), .QN());
   DFF_X1 \buffer_reg[2][4][3][5]  (.D(\input_filter[4][3] [5]), .CK(n_54_4), 
      .Q(\buffer[2][4][3] [5]), .QN());
   DFF_X1 \buffer_reg[2][4][3][4]  (.D(\input_filter[4][3] [4]), .CK(n_54_4), 
      .Q(\buffer[2][4][3] [4]), .QN());
   DFF_X1 \buffer_reg[2][4][3][3]  (.D(\input_filter[4][3] [3]), .CK(n_54_4), 
      .Q(\buffer[2][4][3] [3]), .QN());
   DFF_X1 \buffer_reg[2][4][3][2]  (.D(\input_filter[4][3] [2]), .CK(n_54_4), 
      .Q(\buffer[2][4][3] [2]), .QN());
   DFF_X1 \buffer_reg[2][4][3][1]  (.D(\input_filter[4][3] [1]), .CK(n_54_4), 
      .Q(\buffer[2][4][3] [1]), .QN());
   DFF_X1 \buffer_reg[2][4][3][0]  (.D(\input_filter[4][3] [0]), .CK(n_54_4), 
      .Q(\buffer[2][4][3] [0]), .QN());
   DFF_X1 \buffer_reg[3][4][3][15]  (.D(\input_filter[4][3] [15]), .CK(n_54_5), 
      .Q(\buffer[3][4][3] [15]), .QN());
   DFF_X1 \buffer_reg[3][4][3][14]  (.D(\input_filter[4][3] [14]), .CK(n_54_5), 
      .Q(\buffer[3][4][3] [14]), .QN());
   DFF_X1 \buffer_reg[3][4][3][13]  (.D(\input_filter[4][3] [13]), .CK(n_54_5), 
      .Q(\buffer[3][4][3] [13]), .QN());
   DFF_X1 \buffer_reg[3][4][3][12]  (.D(\input_filter[4][3] [12]), .CK(n_54_5), 
      .Q(\buffer[3][4][3] [12]), .QN());
   DFF_X1 \buffer_reg[3][4][3][11]  (.D(\input_filter[4][3] [11]), .CK(n_54_5), 
      .Q(\buffer[3][4][3] [11]), .QN());
   DFF_X1 \buffer_reg[3][4][3][10]  (.D(\input_filter[4][3] [10]), .CK(n_54_5), 
      .Q(\buffer[3][4][3] [10]), .QN());
   DFF_X1 \buffer_reg[3][4][3][9]  (.D(\input_filter[4][3] [9]), .CK(n_54_5), 
      .Q(\buffer[3][4][3] [9]), .QN());
   DFF_X1 \buffer_reg[3][4][3][8]  (.D(\input_filter[4][3] [8]), .CK(n_54_5), 
      .Q(\buffer[3][4][3] [8]), .QN());
   DFF_X1 \buffer_reg[3][4][3][7]  (.D(\input_filter[4][3] [7]), .CK(n_54_5), 
      .Q(\buffer[3][4][3] [7]), .QN());
   DFF_X1 \buffer_reg[3][4][3][6]  (.D(\input_filter[4][3] [6]), .CK(n_54_5), 
      .Q(\buffer[3][4][3] [6]), .QN());
   DFF_X1 \buffer_reg[3][4][3][5]  (.D(\input_filter[4][3] [5]), .CK(n_54_5), 
      .Q(\buffer[3][4][3] [5]), .QN());
   DFF_X1 \buffer_reg[3][4][3][4]  (.D(\input_filter[4][3] [4]), .CK(n_54_5), 
      .Q(\buffer[3][4][3] [4]), .QN());
   DFF_X1 \buffer_reg[3][4][3][3]  (.D(\input_filter[4][3] [3]), .CK(n_54_5), 
      .Q(\buffer[3][4][3] [3]), .QN());
   DFF_X1 \buffer_reg[3][4][3][2]  (.D(\input_filter[4][3] [2]), .CK(n_54_5), 
      .Q(\buffer[3][4][3] [2]), .QN());
   DFF_X1 \buffer_reg[3][4][3][1]  (.D(\input_filter[4][3] [1]), .CK(n_54_5), 
      .Q(\buffer[3][4][3] [1]), .QN());
   DFF_X1 \buffer_reg[3][4][3][0]  (.D(\input_filter[4][3] [0]), .CK(n_54_5), 
      .Q(\buffer[3][4][3] [0]), .QN());
   DFF_X1 \buffer_reg[13][4][3][15]  (.D(\input_filter[4][3] [15]), .CK(n_54_7), 
      .Q(\buffer[13][4][3] [15]), .QN());
   DFF_X1 \buffer_reg[13][4][3][14]  (.D(\input_filter[4][3] [14]), .CK(n_54_7), 
      .Q(\buffer[13][4][3] [14]), .QN());
   DFF_X1 \buffer_reg[13][4][3][13]  (.D(\input_filter[4][3] [13]), .CK(n_54_7), 
      .Q(\buffer[13][4][3] [13]), .QN());
   DFF_X1 \buffer_reg[13][4][3][12]  (.D(\input_filter[4][3] [12]), .CK(n_54_7), 
      .Q(\buffer[13][4][3] [12]), .QN());
   DFF_X1 \buffer_reg[13][4][3][11]  (.D(\input_filter[4][3] [11]), .CK(n_54_7), 
      .Q(\buffer[13][4][3] [11]), .QN());
   DFF_X1 \buffer_reg[13][4][3][10]  (.D(\input_filter[4][3] [10]), .CK(n_54_7), 
      .Q(\buffer[13][4][3] [10]), .QN());
   DFF_X1 \buffer_reg[13][4][3][9]  (.D(\input_filter[4][3] [9]), .CK(n_54_7), 
      .Q(\buffer[13][4][3] [9]), .QN());
   DFF_X1 \buffer_reg[13][4][3][8]  (.D(\input_filter[4][3] [8]), .CK(n_54_7), 
      .Q(\buffer[13][4][3] [8]), .QN());
   DFF_X1 \buffer_reg[13][4][3][7]  (.D(\input_filter[4][3] [7]), .CK(n_54_7), 
      .Q(\buffer[13][4][3] [7]), .QN());
   DFF_X1 \buffer_reg[13][4][3][6]  (.D(\input_filter[4][3] [6]), .CK(n_54_7), 
      .Q(\buffer[13][4][3] [6]), .QN());
   DFF_X1 \buffer_reg[13][4][3][5]  (.D(\input_filter[4][3] [5]), .CK(n_54_7), 
      .Q(\buffer[13][4][3] [5]), .QN());
   DFF_X1 \buffer_reg[13][4][3][4]  (.D(\input_filter[4][3] [4]), .CK(n_54_7), 
      .Q(\buffer[13][4][3] [4]), .QN());
   DFF_X1 \buffer_reg[13][4][3][3]  (.D(\input_filter[4][3] [3]), .CK(n_54_7), 
      .Q(\buffer[13][4][3] [3]), .QN());
   DFF_X1 \buffer_reg[13][4][3][2]  (.D(\input_filter[4][3] [2]), .CK(n_54_7), 
      .Q(\buffer[13][4][3] [2]), .QN());
   DFF_X1 \buffer_reg[13][4][3][1]  (.D(\input_filter[4][3] [1]), .CK(n_54_7), 
      .Q(\buffer[13][4][3] [1]), .QN());
   DFF_X1 \buffer_reg[13][4][3][0]  (.D(\input_filter[4][3] [0]), .CK(n_54_7), 
      .Q(\buffer[13][4][3] [0]), .QN());
   DFF_X1 \buffer_reg[14][4][3][15]  (.D(\input_filter[4][3] [15]), .CK(n_54_8), 
      .Q(\buffer[14][4][3] [15]), .QN());
   DFF_X1 \buffer_reg[14][4][3][14]  (.D(\input_filter[4][3] [14]), .CK(n_54_8), 
      .Q(\buffer[14][4][3] [14]), .QN());
   DFF_X1 \buffer_reg[14][4][3][13]  (.D(\input_filter[4][3] [13]), .CK(n_54_8), 
      .Q(\buffer[14][4][3] [13]), .QN());
   DFF_X1 \buffer_reg[14][4][3][12]  (.D(\input_filter[4][3] [12]), .CK(n_54_8), 
      .Q(\buffer[14][4][3] [12]), .QN());
   DFF_X1 \buffer_reg[14][4][3][11]  (.D(\input_filter[4][3] [11]), .CK(n_54_8), 
      .Q(\buffer[14][4][3] [11]), .QN());
   DFF_X1 \buffer_reg[14][4][3][10]  (.D(\input_filter[4][3] [10]), .CK(n_54_8), 
      .Q(\buffer[14][4][3] [10]), .QN());
   DFF_X1 \buffer_reg[14][4][3][9]  (.D(\input_filter[4][3] [9]), .CK(n_54_8), 
      .Q(\buffer[14][4][3] [9]), .QN());
   DFF_X1 \buffer_reg[14][4][3][8]  (.D(\input_filter[4][3] [8]), .CK(n_54_8), 
      .Q(\buffer[14][4][3] [8]), .QN());
   DFF_X1 \buffer_reg[14][4][3][7]  (.D(\input_filter[4][3] [7]), .CK(n_54_8), 
      .Q(\buffer[14][4][3] [7]), .QN());
   DFF_X1 \buffer_reg[14][4][3][6]  (.D(\input_filter[4][3] [6]), .CK(n_54_8), 
      .Q(\buffer[14][4][3] [6]), .QN());
   DFF_X1 \buffer_reg[14][4][3][5]  (.D(\input_filter[4][3] [5]), .CK(n_54_8), 
      .Q(\buffer[14][4][3] [5]), .QN());
   DFF_X1 \buffer_reg[14][4][3][4]  (.D(\input_filter[4][3] [4]), .CK(n_54_8), 
      .Q(\buffer[14][4][3] [4]), .QN());
   DFF_X1 \buffer_reg[14][4][3][3]  (.D(\input_filter[4][3] [3]), .CK(n_54_8), 
      .Q(\buffer[14][4][3] [3]), .QN());
   DFF_X1 \buffer_reg[14][4][3][2]  (.D(\input_filter[4][3] [2]), .CK(n_54_8), 
      .Q(\buffer[14][4][3] [2]), .QN());
   DFF_X1 \buffer_reg[14][4][3][1]  (.D(\input_filter[4][3] [1]), .CK(n_54_8), 
      .Q(\buffer[14][4][3] [1]), .QN());
   DFF_X1 \buffer_reg[14][4][3][0]  (.D(\input_filter[4][3] [0]), .CK(n_54_8), 
      .Q(\buffer[14][4][3] [0]), .QN());
   DFF_X1 \buffer_reg[15][4][3][15]  (.D(\input_filter[4][3] [15]), .CK(n_54_9), 
      .Q(\buffer[15][4][3] [15]), .QN());
   DFF_X1 \buffer_reg[15][4][3][14]  (.D(\input_filter[4][3] [14]), .CK(n_54_9), 
      .Q(\buffer[15][4][3] [14]), .QN());
   DFF_X1 \buffer_reg[15][4][3][13]  (.D(\input_filter[4][3] [13]), .CK(n_54_9), 
      .Q(\buffer[15][4][3] [13]), .QN());
   DFF_X1 \buffer_reg[15][4][3][12]  (.D(\input_filter[4][3] [12]), .CK(n_54_9), 
      .Q(\buffer[15][4][3] [12]), .QN());
   DFF_X1 \buffer_reg[15][4][3][11]  (.D(\input_filter[4][3] [11]), .CK(n_54_9), 
      .Q(\buffer[15][4][3] [11]), .QN());
   DFF_X1 \buffer_reg[15][4][3][10]  (.D(\input_filter[4][3] [10]), .CK(n_54_9), 
      .Q(\buffer[15][4][3] [10]), .QN());
   DFF_X1 \buffer_reg[15][4][3][9]  (.D(\input_filter[4][3] [9]), .CK(n_54_9), 
      .Q(\buffer[15][4][3] [9]), .QN());
   DFF_X1 \buffer_reg[15][4][3][8]  (.D(\input_filter[4][3] [8]), .CK(n_54_9), 
      .Q(\buffer[15][4][3] [8]), .QN());
   DFF_X1 \buffer_reg[15][4][3][7]  (.D(\input_filter[4][3] [7]), .CK(n_54_9), 
      .Q(\buffer[15][4][3] [7]), .QN());
   DFF_X1 \buffer_reg[15][4][3][6]  (.D(\input_filter[4][3] [6]), .CK(n_54_9), 
      .Q(\buffer[15][4][3] [6]), .QN());
   DFF_X1 \buffer_reg[15][4][3][5]  (.D(\input_filter[4][3] [5]), .CK(n_54_9), 
      .Q(\buffer[15][4][3] [5]), .QN());
   DFF_X1 \buffer_reg[15][4][3][4]  (.D(\input_filter[4][3] [4]), .CK(n_54_9), 
      .Q(\buffer[15][4][3] [4]), .QN());
   DFF_X1 \buffer_reg[15][4][3][3]  (.D(\input_filter[4][3] [3]), .CK(n_54_9), 
      .Q(\buffer[15][4][3] [3]), .QN());
   DFF_X1 \buffer_reg[15][4][3][2]  (.D(\input_filter[4][3] [2]), .CK(n_54_9), 
      .Q(\buffer[15][4][3] [2]), .QN());
   DFF_X1 \buffer_reg[15][4][3][1]  (.D(\input_filter[4][3] [1]), .CK(n_54_9), 
      .Q(\buffer[15][4][3] [1]), .QN());
   DFF_X1 \buffer_reg[15][4][3][0]  (.D(\input_filter[4][3] [0]), .CK(n_54_9), 
      .Q(\buffer[15][4][3] [0]), .QN());
   CLKGATETST_X1 \clk_gate_buffer_reg[0][4][4]_reg  (.CK(read), .E(n_0), 
      .SE(1'b0), .GCK(n_54_6));
   DFF_X1 \buffer_reg[0][4][4][15]  (.D(\input_filter[4][4] [15]), .CK(n_54_6), 
      .Q(\buffer[0][4][4] [15]), .QN());
   DFF_X1 \buffer_reg[0][4][4][14]  (.D(\input_filter[4][4] [14]), .CK(n_54_6), 
      .Q(\buffer[0][4][4] [14]), .QN());
   DFF_X1 \buffer_reg[0][4][4][13]  (.D(\input_filter[4][4] [13]), .CK(n_54_6), 
      .Q(\buffer[0][4][4] [13]), .QN());
   DFF_X1 \buffer_reg[0][4][4][12]  (.D(\input_filter[4][4] [12]), .CK(n_54_6), 
      .Q(\buffer[0][4][4] [12]), .QN());
   DFF_X1 \buffer_reg[0][4][4][11]  (.D(\input_filter[4][4] [11]), .CK(n_54_6), 
      .Q(\buffer[0][4][4] [11]), .QN());
   DFF_X1 \buffer_reg[0][4][4][10]  (.D(\input_filter[4][4] [10]), .CK(n_54_6), 
      .Q(\buffer[0][4][4] [10]), .QN());
   DFF_X1 \buffer_reg[0][4][4][9]  (.D(\input_filter[4][4] [9]), .CK(n_54_6), 
      .Q(\buffer[0][4][4] [9]), .QN());
   DFF_X1 \buffer_reg[0][4][4][8]  (.D(\input_filter[4][4] [8]), .CK(n_54_6), 
      .Q(\buffer[0][4][4] [8]), .QN());
   DFF_X1 \buffer_reg[0][4][4][7]  (.D(\input_filter[4][4] [7]), .CK(n_54_6), 
      .Q(\buffer[0][4][4] [7]), .QN());
   DFF_X1 \buffer_reg[0][4][4][6]  (.D(\input_filter[4][4] [6]), .CK(n_54_6), 
      .Q(\buffer[0][4][4] [6]), .QN());
   DFF_X1 \buffer_reg[0][4][4][5]  (.D(\input_filter[4][4] [5]), .CK(n_54_6), 
      .Q(\buffer[0][4][4] [5]), .QN());
   DFF_X1 \buffer_reg[0][4][4][4]  (.D(\input_filter[4][4] [4]), .CK(n_54_6), 
      .Q(\buffer[0][4][4] [4]), .QN());
   DFF_X1 \buffer_reg[0][4][4][3]  (.D(\input_filter[4][4] [3]), .CK(n_54_6), 
      .Q(\buffer[0][4][4] [3]), .QN());
   DFF_X1 \buffer_reg[0][4][4][2]  (.D(\input_filter[4][4] [2]), .CK(n_54_6), 
      .Q(\buffer[0][4][4] [2]), .QN());
   DFF_X1 \buffer_reg[0][4][4][1]  (.D(\input_filter[4][4] [1]), .CK(n_54_6), 
      .Q(\buffer[0][4][4] [1]), .QN());
   DFF_X1 \buffer_reg[0][4][4][0]  (.D(\input_filter[4][4] [0]), .CK(n_54_6), 
      .Q(\buffer[0][4][4] [0]), .QN());
   DFF_X1 \buffer_reg[1][4][4][15]  (.D(\input_filter[4][4] [15]), .CK(n_54_3), 
      .Q(\buffer[1][4][4] [15]), .QN());
   DFF_X1 \buffer_reg[1][4][4][14]  (.D(\input_filter[4][4] [14]), .CK(n_54_3), 
      .Q(\buffer[1][4][4] [14]), .QN());
   DFF_X1 \buffer_reg[1][4][4][13]  (.D(\input_filter[4][4] [13]), .CK(n_54_3), 
      .Q(\buffer[1][4][4] [13]), .QN());
   DFF_X1 \buffer_reg[1][4][4][12]  (.D(\input_filter[4][4] [12]), .CK(n_54_3), 
      .Q(\buffer[1][4][4] [12]), .QN());
   DFF_X1 \buffer_reg[1][4][4][11]  (.D(\input_filter[4][4] [11]), .CK(n_54_3), 
      .Q(\buffer[1][4][4] [11]), .QN());
   DFF_X1 \buffer_reg[1][4][4][10]  (.D(\input_filter[4][4] [10]), .CK(n_54_3), 
      .Q(\buffer[1][4][4] [10]), .QN());
   DFF_X1 \buffer_reg[1][4][4][9]  (.D(\input_filter[4][4] [9]), .CK(n_54_3), 
      .Q(\buffer[1][4][4] [9]), .QN());
   DFF_X1 \buffer_reg[1][4][4][8]  (.D(\input_filter[4][4] [8]), .CK(n_54_3), 
      .Q(\buffer[1][4][4] [8]), .QN());
   DFF_X1 \buffer_reg[1][4][4][7]  (.D(\input_filter[4][4] [7]), .CK(n_54_3), 
      .Q(\buffer[1][4][4] [7]), .QN());
   DFF_X1 \buffer_reg[1][4][4][6]  (.D(\input_filter[4][4] [6]), .CK(n_54_3), 
      .Q(\buffer[1][4][4] [6]), .QN());
   DFF_X1 \buffer_reg[1][4][4][5]  (.D(\input_filter[4][4] [5]), .CK(n_54_3), 
      .Q(\buffer[1][4][4] [5]), .QN());
   DFF_X1 \buffer_reg[1][4][4][4]  (.D(\input_filter[4][4] [4]), .CK(n_54_3), 
      .Q(\buffer[1][4][4] [4]), .QN());
   DFF_X1 \buffer_reg[1][4][4][3]  (.D(\input_filter[4][4] [3]), .CK(n_54_3), 
      .Q(\buffer[1][4][4] [3]), .QN());
   DFF_X1 \buffer_reg[1][4][4][2]  (.D(\input_filter[4][4] [2]), .CK(n_54_3), 
      .Q(\buffer[1][4][4] [2]), .QN());
   DFF_X1 \buffer_reg[1][4][4][1]  (.D(\input_filter[4][4] [1]), .CK(n_54_3), 
      .Q(\buffer[1][4][4] [1]), .QN());
   DFF_X1 \buffer_reg[1][4][4][0]  (.D(\input_filter[4][4] [0]), .CK(n_54_3), 
      .Q(\buffer[1][4][4] [0]), .QN());
   DFF_X1 \buffer_reg[2][4][4][15]  (.D(\input_filter[4][4] [15]), .CK(n_54_4), 
      .Q(\buffer[2][4][4] [15]), .QN());
   DFF_X1 \buffer_reg[2][4][4][14]  (.D(\input_filter[4][4] [14]), .CK(n_54_4), 
      .Q(\buffer[2][4][4] [14]), .QN());
   DFF_X1 \buffer_reg[2][4][4][13]  (.D(\input_filter[4][4] [13]), .CK(n_54_4), 
      .Q(\buffer[2][4][4] [13]), .QN());
   DFF_X1 \buffer_reg[2][4][4][12]  (.D(\input_filter[4][4] [12]), .CK(n_54_4), 
      .Q(\buffer[2][4][4] [12]), .QN());
   DFF_X1 \buffer_reg[2][4][4][11]  (.D(\input_filter[4][4] [11]), .CK(n_54_4), 
      .Q(\buffer[2][4][4] [11]), .QN());
   DFF_X1 \buffer_reg[2][4][4][10]  (.D(\input_filter[4][4] [10]), .CK(n_54_4), 
      .Q(\buffer[2][4][4] [10]), .QN());
   DFF_X1 \buffer_reg[2][4][4][9]  (.D(\input_filter[4][4] [9]), .CK(n_54_4), 
      .Q(\buffer[2][4][4] [9]), .QN());
   DFF_X1 \buffer_reg[2][4][4][8]  (.D(\input_filter[4][4] [8]), .CK(n_54_4), 
      .Q(\buffer[2][4][4] [8]), .QN());
   DFF_X1 \buffer_reg[2][4][4][7]  (.D(\input_filter[4][4] [7]), .CK(n_54_4), 
      .Q(\buffer[2][4][4] [7]), .QN());
   DFF_X1 \buffer_reg[2][4][4][6]  (.D(\input_filter[4][4] [6]), .CK(n_54_4), 
      .Q(\buffer[2][4][4] [6]), .QN());
   DFF_X1 \buffer_reg[2][4][4][5]  (.D(\input_filter[4][4] [5]), .CK(n_54_4), 
      .Q(\buffer[2][4][4] [5]), .QN());
   DFF_X1 \buffer_reg[2][4][4][4]  (.D(\input_filter[4][4] [4]), .CK(n_54_4), 
      .Q(\buffer[2][4][4] [4]), .QN());
   DFF_X1 \buffer_reg[2][4][4][3]  (.D(\input_filter[4][4] [3]), .CK(n_54_4), 
      .Q(\buffer[2][4][4] [3]), .QN());
   DFF_X1 \buffer_reg[2][4][4][2]  (.D(\input_filter[4][4] [2]), .CK(n_54_4), 
      .Q(\buffer[2][4][4] [2]), .QN());
   DFF_X1 \buffer_reg[2][4][4][1]  (.D(\input_filter[4][4] [1]), .CK(n_54_4), 
      .Q(\buffer[2][4][4] [1]), .QN());
   DFF_X1 \buffer_reg[2][4][4][0]  (.D(\input_filter[4][4] [0]), .CK(n_54_4), 
      .Q(\buffer[2][4][4] [0]), .QN());
   DFF_X1 \buffer_reg[3][4][4][15]  (.D(\input_filter[4][4] [15]), .CK(n_54_5), 
      .Q(\buffer[3][4][4] [15]), .QN());
   DFF_X1 \buffer_reg[3][4][4][14]  (.D(\input_filter[4][4] [14]), .CK(n_54_5), 
      .Q(\buffer[3][4][4] [14]), .QN());
   DFF_X1 \buffer_reg[3][4][4][13]  (.D(\input_filter[4][4] [13]), .CK(n_54_5), 
      .Q(\buffer[3][4][4] [13]), .QN());
   DFF_X1 \buffer_reg[3][4][4][12]  (.D(\input_filter[4][4] [12]), .CK(n_54_5), 
      .Q(\buffer[3][4][4] [12]), .QN());
   DFF_X1 \buffer_reg[3][4][4][11]  (.D(\input_filter[4][4] [11]), .CK(n_54_5), 
      .Q(\buffer[3][4][4] [11]), .QN());
   DFF_X1 \buffer_reg[3][4][4][10]  (.D(\input_filter[4][4] [10]), .CK(n_54_5), 
      .Q(\buffer[3][4][4] [10]), .QN());
   DFF_X1 \buffer_reg[3][4][4][9]  (.D(\input_filter[4][4] [9]), .CK(n_54_5), 
      .Q(\buffer[3][4][4] [9]), .QN());
   DFF_X1 \buffer_reg[3][4][4][8]  (.D(\input_filter[4][4] [8]), .CK(n_54_5), 
      .Q(\buffer[3][4][4] [8]), .QN());
   DFF_X1 \buffer_reg[3][4][4][7]  (.D(\input_filter[4][4] [7]), .CK(n_54_5), 
      .Q(\buffer[3][4][4] [7]), .QN());
   DFF_X1 \buffer_reg[3][4][4][6]  (.D(\input_filter[4][4] [6]), .CK(n_54_5), 
      .Q(\buffer[3][4][4] [6]), .QN());
   DFF_X1 \buffer_reg[3][4][4][5]  (.D(\input_filter[4][4] [5]), .CK(n_54_5), 
      .Q(\buffer[3][4][4] [5]), .QN());
   DFF_X1 \buffer_reg[3][4][4][4]  (.D(\input_filter[4][4] [4]), .CK(n_54_5), 
      .Q(\buffer[3][4][4] [4]), .QN());
   DFF_X1 \buffer_reg[3][4][4][3]  (.D(\input_filter[4][4] [3]), .CK(n_54_5), 
      .Q(\buffer[3][4][4] [3]), .QN());
   DFF_X1 \buffer_reg[3][4][4][2]  (.D(\input_filter[4][4] [2]), .CK(n_54_5), 
      .Q(\buffer[3][4][4] [2]), .QN());
   DFF_X1 \buffer_reg[3][4][4][1]  (.D(\input_filter[4][4] [1]), .CK(n_54_5), 
      .Q(\buffer[3][4][4] [1]), .QN());
   DFF_X1 \buffer_reg[3][4][4][0]  (.D(\input_filter[4][4] [0]), .CK(n_54_5), 
      .Q(\buffer[3][4][4] [0]), .QN());
   CLKGATETST_X1 \clk_gate_buffer_reg[4][4][4]_reg  (.CK(read), .E(n_4), 
      .SE(1'b0), .GCK(n_54_10));
   DFF_X1 \buffer_reg[4][4][4][15]  (.D(\input_filter[4][4] [15]), .CK(n_54_10), 
      .Q(\buffer[4][4][4] [15]), .QN());
   DFF_X1 \buffer_reg[4][4][4][14]  (.D(\input_filter[4][4] [14]), .CK(n_54_10), 
      .Q(\buffer[4][4][4] [14]), .QN());
   DFF_X1 \buffer_reg[4][4][4][13]  (.D(\input_filter[4][4] [13]), .CK(n_54_10), 
      .Q(\buffer[4][4][4] [13]), .QN());
   DFF_X1 \buffer_reg[4][4][4][12]  (.D(\input_filter[4][4] [12]), .CK(n_54_10), 
      .Q(\buffer[4][4][4] [12]), .QN());
   DFF_X1 \buffer_reg[4][4][4][11]  (.D(\input_filter[4][4] [11]), .CK(n_54_10), 
      .Q(\buffer[4][4][4] [11]), .QN());
   DFF_X1 \buffer_reg[4][4][4][10]  (.D(\input_filter[4][4] [10]), .CK(n_54_10), 
      .Q(\buffer[4][4][4] [10]), .QN());
   DFF_X1 \buffer_reg[4][4][4][9]  (.D(\input_filter[4][4] [9]), .CK(n_54_10), 
      .Q(\buffer[4][4][4] [9]), .QN());
   DFF_X1 \buffer_reg[4][4][4][8]  (.D(\input_filter[4][4] [8]), .CK(n_54_10), 
      .Q(\buffer[4][4][4] [8]), .QN());
   DFF_X1 \buffer_reg[4][4][4][7]  (.D(\input_filter[4][4] [7]), .CK(n_54_10), 
      .Q(\buffer[4][4][4] [7]), .QN());
   DFF_X1 \buffer_reg[4][4][4][6]  (.D(\input_filter[4][4] [6]), .CK(n_54_10), 
      .Q(\buffer[4][4][4] [6]), .QN());
   DFF_X1 \buffer_reg[4][4][4][5]  (.D(\input_filter[4][4] [5]), .CK(n_54_10), 
      .Q(\buffer[4][4][4] [5]), .QN());
   DFF_X1 \buffer_reg[4][4][4][4]  (.D(\input_filter[4][4] [4]), .CK(n_54_10), 
      .Q(\buffer[4][4][4] [4]), .QN());
   DFF_X1 \buffer_reg[4][4][4][3]  (.D(\input_filter[4][4] [3]), .CK(n_54_10), 
      .Q(\buffer[4][4][4] [3]), .QN());
   DFF_X1 \buffer_reg[4][4][4][2]  (.D(\input_filter[4][4] [2]), .CK(n_54_10), 
      .Q(\buffer[4][4][4] [2]), .QN());
   DFF_X1 \buffer_reg[4][4][4][1]  (.D(\input_filter[4][4] [1]), .CK(n_54_10), 
      .Q(\buffer[4][4][4] [1]), .QN());
   DFF_X1 \buffer_reg[4][4][4][0]  (.D(\input_filter[4][4] [0]), .CK(n_54_10), 
      .Q(\buffer[4][4][4] [0]), .QN());
   CLKGATETST_X1 \clk_gate_buffer_reg[5][4][4]_reg  (.CK(read), .E(n_5), 
      .SE(1'b0), .GCK(n_54_11));
   DFF_X1 \buffer_reg[5][4][4][15]  (.D(\input_filter[4][4] [15]), .CK(n_54_11), 
      .Q(\buffer[5][4][4] [15]), .QN());
   DFF_X1 \buffer_reg[5][4][4][14]  (.D(\input_filter[4][4] [14]), .CK(n_54_11), 
      .Q(\buffer[5][4][4] [14]), .QN());
   DFF_X1 \buffer_reg[5][4][4][13]  (.D(\input_filter[4][4] [13]), .CK(n_54_11), 
      .Q(\buffer[5][4][4] [13]), .QN());
   DFF_X1 \buffer_reg[5][4][4][12]  (.D(\input_filter[4][4] [12]), .CK(n_54_11), 
      .Q(\buffer[5][4][4] [12]), .QN());
   DFF_X1 \buffer_reg[5][4][4][11]  (.D(\input_filter[4][4] [11]), .CK(n_54_11), 
      .Q(\buffer[5][4][4] [11]), .QN());
   DFF_X1 \buffer_reg[5][4][4][10]  (.D(\input_filter[4][4] [10]), .CK(n_54_11), 
      .Q(\buffer[5][4][4] [10]), .QN());
   DFF_X1 \buffer_reg[5][4][4][9]  (.D(\input_filter[4][4] [9]), .CK(n_54_11), 
      .Q(\buffer[5][4][4] [9]), .QN());
   DFF_X1 \buffer_reg[5][4][4][8]  (.D(\input_filter[4][4] [8]), .CK(n_54_11), 
      .Q(\buffer[5][4][4] [8]), .QN());
   DFF_X1 \buffer_reg[5][4][4][7]  (.D(\input_filter[4][4] [7]), .CK(n_54_11), 
      .Q(\buffer[5][4][4] [7]), .QN());
   DFF_X1 \buffer_reg[5][4][4][6]  (.D(\input_filter[4][4] [6]), .CK(n_54_11), 
      .Q(\buffer[5][4][4] [6]), .QN());
   DFF_X1 \buffer_reg[5][4][4][5]  (.D(\input_filter[4][4] [5]), .CK(n_54_11), 
      .Q(\buffer[5][4][4] [5]), .QN());
   DFF_X1 \buffer_reg[5][4][4][4]  (.D(\input_filter[4][4] [4]), .CK(n_54_11), 
      .Q(\buffer[5][4][4] [4]), .QN());
   DFF_X1 \buffer_reg[5][4][4][3]  (.D(\input_filter[4][4] [3]), .CK(n_54_11), 
      .Q(\buffer[5][4][4] [3]), .QN());
   DFF_X1 \buffer_reg[5][4][4][2]  (.D(\input_filter[4][4] [2]), .CK(n_54_11), 
      .Q(\buffer[5][4][4] [2]), .QN());
   DFF_X1 \buffer_reg[5][4][4][1]  (.D(\input_filter[4][4] [1]), .CK(n_54_11), 
      .Q(\buffer[5][4][4] [1]), .QN());
   DFF_X1 \buffer_reg[5][4][4][0]  (.D(\input_filter[4][4] [0]), .CK(n_54_11), 
      .Q(\buffer[5][4][4] [0]), .QN());
   CLKGATETST_X1 \clk_gate_buffer_reg[6][4][4]_reg  (.CK(read), .E(n_6), 
      .SE(1'b0), .GCK(n_54_12));
   DFF_X1 \buffer_reg[6][4][4][15]  (.D(\input_filter[4][4] [15]), .CK(n_54_12), 
      .Q(\buffer[6][4][4] [15]), .QN());
   DFF_X1 \buffer_reg[6][4][4][14]  (.D(\input_filter[4][4] [14]), .CK(n_54_12), 
      .Q(\buffer[6][4][4] [14]), .QN());
   DFF_X1 \buffer_reg[6][4][4][13]  (.D(\input_filter[4][4] [13]), .CK(n_54_12), 
      .Q(\buffer[6][4][4] [13]), .QN());
   DFF_X1 \buffer_reg[6][4][4][12]  (.D(\input_filter[4][4] [12]), .CK(n_54_12), 
      .Q(\buffer[6][4][4] [12]), .QN());
   DFF_X1 \buffer_reg[6][4][4][11]  (.D(\input_filter[4][4] [11]), .CK(n_54_12), 
      .Q(\buffer[6][4][4] [11]), .QN());
   DFF_X1 \buffer_reg[6][4][4][10]  (.D(\input_filter[4][4] [10]), .CK(n_54_12), 
      .Q(\buffer[6][4][4] [10]), .QN());
   DFF_X1 \buffer_reg[6][4][4][9]  (.D(\input_filter[4][4] [9]), .CK(n_54_12), 
      .Q(\buffer[6][4][4] [9]), .QN());
   DFF_X1 \buffer_reg[6][4][4][8]  (.D(\input_filter[4][4] [8]), .CK(n_54_12), 
      .Q(\buffer[6][4][4] [8]), .QN());
   DFF_X1 \buffer_reg[6][4][4][7]  (.D(\input_filter[4][4] [7]), .CK(n_54_12), 
      .Q(\buffer[6][4][4] [7]), .QN());
   DFF_X1 \buffer_reg[6][4][4][6]  (.D(\input_filter[4][4] [6]), .CK(n_54_12), 
      .Q(\buffer[6][4][4] [6]), .QN());
   DFF_X1 \buffer_reg[6][4][4][5]  (.D(\input_filter[4][4] [5]), .CK(n_54_12), 
      .Q(\buffer[6][4][4] [5]), .QN());
   DFF_X1 \buffer_reg[6][4][4][4]  (.D(\input_filter[4][4] [4]), .CK(n_54_12), 
      .Q(\buffer[6][4][4] [4]), .QN());
   DFF_X1 \buffer_reg[6][4][4][3]  (.D(\input_filter[4][4] [3]), .CK(n_54_12), 
      .Q(\buffer[6][4][4] [3]), .QN());
   DFF_X1 \buffer_reg[6][4][4][2]  (.D(\input_filter[4][4] [2]), .CK(n_54_12), 
      .Q(\buffer[6][4][4] [2]), .QN());
   DFF_X1 \buffer_reg[6][4][4][1]  (.D(\input_filter[4][4] [1]), .CK(n_54_12), 
      .Q(\buffer[6][4][4] [1]), .QN());
   DFF_X1 \buffer_reg[6][4][4][0]  (.D(\input_filter[4][4] [0]), .CK(n_54_12), 
      .Q(\buffer[6][4][4] [0]), .QN());
   CLKGATETST_X1 \clk_gate_buffer_reg[7][4][4]_reg  (.CK(read), .E(n_7), 
      .SE(1'b0), .GCK(n_54_13));
   DFF_X1 \buffer_reg[7][4][4][15]  (.D(\input_filter[4][4] [15]), .CK(n_54_13), 
      .Q(\buffer[7][4][4] [15]), .QN());
   DFF_X1 \buffer_reg[7][4][4][14]  (.D(\input_filter[4][4] [14]), .CK(n_54_13), 
      .Q(\buffer[7][4][4] [14]), .QN());
   DFF_X1 \buffer_reg[7][4][4][13]  (.D(\input_filter[4][4] [13]), .CK(n_54_13), 
      .Q(\buffer[7][4][4] [13]), .QN());
   DFF_X1 \buffer_reg[7][4][4][12]  (.D(\input_filter[4][4] [12]), .CK(n_54_13), 
      .Q(\buffer[7][4][4] [12]), .QN());
   DFF_X1 \buffer_reg[7][4][4][11]  (.D(\input_filter[4][4] [11]), .CK(n_54_13), 
      .Q(\buffer[7][4][4] [11]), .QN());
   DFF_X1 \buffer_reg[7][4][4][10]  (.D(\input_filter[4][4] [10]), .CK(n_54_13), 
      .Q(\buffer[7][4][4] [10]), .QN());
   DFF_X1 \buffer_reg[7][4][4][9]  (.D(\input_filter[4][4] [9]), .CK(n_54_13), 
      .Q(\buffer[7][4][4] [9]), .QN());
   DFF_X1 \buffer_reg[7][4][4][8]  (.D(\input_filter[4][4] [8]), .CK(n_54_13), 
      .Q(\buffer[7][4][4] [8]), .QN());
   DFF_X1 \buffer_reg[7][4][4][7]  (.D(\input_filter[4][4] [7]), .CK(n_54_13), 
      .Q(\buffer[7][4][4] [7]), .QN());
   DFF_X1 \buffer_reg[7][4][4][6]  (.D(\input_filter[4][4] [6]), .CK(n_54_13), 
      .Q(\buffer[7][4][4] [6]), .QN());
   DFF_X1 \buffer_reg[7][4][4][5]  (.D(\input_filter[4][4] [5]), .CK(n_54_13), 
      .Q(\buffer[7][4][4] [5]), .QN());
   DFF_X1 \buffer_reg[7][4][4][4]  (.D(\input_filter[4][4] [4]), .CK(n_54_13), 
      .Q(\buffer[7][4][4] [4]), .QN());
   DFF_X1 \buffer_reg[7][4][4][3]  (.D(\input_filter[4][4] [3]), .CK(n_54_13), 
      .Q(\buffer[7][4][4] [3]), .QN());
   DFF_X1 \buffer_reg[7][4][4][2]  (.D(\input_filter[4][4] [2]), .CK(n_54_13), 
      .Q(\buffer[7][4][4] [2]), .QN());
   DFF_X1 \buffer_reg[7][4][4][1]  (.D(\input_filter[4][4] [1]), .CK(n_54_13), 
      .Q(\buffer[7][4][4] [1]), .QN());
   DFF_X1 \buffer_reg[7][4][4][0]  (.D(\input_filter[4][4] [0]), .CK(n_54_13), 
      .Q(\buffer[7][4][4] [0]), .QN());
   CLKGATETST_X1 \clk_gate_buffer_reg[8][4][4]_reg  (.CK(read), .E(n_8), 
      .SE(1'b0), .GCK(n_54_14));
   DFF_X1 \buffer_reg[8][4][4][15]  (.D(\input_filter[4][4] [15]), .CK(n_54_14), 
      .Q(\buffer[8][4][4] [15]), .QN());
   DFF_X1 \buffer_reg[8][4][4][14]  (.D(\input_filter[4][4] [14]), .CK(n_54_14), 
      .Q(\buffer[8][4][4] [14]), .QN());
   DFF_X1 \buffer_reg[8][4][4][13]  (.D(\input_filter[4][4] [13]), .CK(n_54_14), 
      .Q(\buffer[8][4][4] [13]), .QN());
   DFF_X1 \buffer_reg[8][4][4][12]  (.D(\input_filter[4][4] [12]), .CK(n_54_14), 
      .Q(\buffer[8][4][4] [12]), .QN());
   DFF_X1 \buffer_reg[8][4][4][11]  (.D(\input_filter[4][4] [11]), .CK(n_54_14), 
      .Q(\buffer[8][4][4] [11]), .QN());
   DFF_X1 \buffer_reg[8][4][4][10]  (.D(\input_filter[4][4] [10]), .CK(n_54_14), 
      .Q(\buffer[8][4][4] [10]), .QN());
   DFF_X1 \buffer_reg[8][4][4][9]  (.D(\input_filter[4][4] [9]), .CK(n_54_14), 
      .Q(\buffer[8][4][4] [9]), .QN());
   DFF_X1 \buffer_reg[8][4][4][8]  (.D(\input_filter[4][4] [8]), .CK(n_54_14), 
      .Q(\buffer[8][4][4] [8]), .QN());
   DFF_X1 \buffer_reg[8][4][4][7]  (.D(\input_filter[4][4] [7]), .CK(n_54_14), 
      .Q(\buffer[8][4][4] [7]), .QN());
   DFF_X1 \buffer_reg[8][4][4][6]  (.D(\input_filter[4][4] [6]), .CK(n_54_14), 
      .Q(\buffer[8][4][4] [6]), .QN());
   DFF_X1 \buffer_reg[8][4][4][5]  (.D(\input_filter[4][4] [5]), .CK(n_54_14), 
      .Q(\buffer[8][4][4] [5]), .QN());
   DFF_X1 \buffer_reg[8][4][4][4]  (.D(\input_filter[4][4] [4]), .CK(n_54_14), 
      .Q(\buffer[8][4][4] [4]), .QN());
   DFF_X1 \buffer_reg[8][4][4][3]  (.D(\input_filter[4][4] [3]), .CK(n_54_14), 
      .Q(\buffer[8][4][4] [3]), .QN());
   DFF_X1 \buffer_reg[8][4][4][2]  (.D(\input_filter[4][4] [2]), .CK(n_54_14), 
      .Q(\buffer[8][4][4] [2]), .QN());
   DFF_X1 \buffer_reg[8][4][4][1]  (.D(\input_filter[4][4] [1]), .CK(n_54_14), 
      .Q(\buffer[8][4][4] [1]), .QN());
   DFF_X1 \buffer_reg[8][4][4][0]  (.D(\input_filter[4][4] [0]), .CK(n_54_14), 
      .Q(\buffer[8][4][4] [0]), .QN());
   CLKGATETST_X1 \clk_gate_buffer_reg[9][4][4]_reg  (.CK(read), .E(n_9), 
      .SE(1'b0), .GCK(n_54_15));
   DFF_X1 \buffer_reg[9][4][4][15]  (.D(\input_filter[4][4] [15]), .CK(n_54_15), 
      .Q(\buffer[9][4][4] [15]), .QN());
   DFF_X1 \buffer_reg[9][4][4][14]  (.D(\input_filter[4][4] [14]), .CK(n_54_15), 
      .Q(\buffer[9][4][4] [14]), .QN());
   DFF_X1 \buffer_reg[9][4][4][13]  (.D(\input_filter[4][4] [13]), .CK(n_54_15), 
      .Q(\buffer[9][4][4] [13]), .QN());
   DFF_X1 \buffer_reg[9][4][4][12]  (.D(\input_filter[4][4] [12]), .CK(n_54_15), 
      .Q(\buffer[9][4][4] [12]), .QN());
   DFF_X1 \buffer_reg[9][4][4][11]  (.D(\input_filter[4][4] [11]), .CK(n_54_15), 
      .Q(\buffer[9][4][4] [11]), .QN());
   DFF_X1 \buffer_reg[9][4][4][10]  (.D(\input_filter[4][4] [10]), .CK(n_54_15), 
      .Q(\buffer[9][4][4] [10]), .QN());
   DFF_X1 \buffer_reg[9][4][4][9]  (.D(\input_filter[4][4] [9]), .CK(n_54_15), 
      .Q(\buffer[9][4][4] [9]), .QN());
   DFF_X1 \buffer_reg[9][4][4][8]  (.D(\input_filter[4][4] [8]), .CK(n_54_15), 
      .Q(\buffer[9][4][4] [8]), .QN());
   DFF_X1 \buffer_reg[9][4][4][7]  (.D(\input_filter[4][4] [7]), .CK(n_54_15), 
      .Q(\buffer[9][4][4] [7]), .QN());
   DFF_X1 \buffer_reg[9][4][4][6]  (.D(\input_filter[4][4] [6]), .CK(n_54_15), 
      .Q(\buffer[9][4][4] [6]), .QN());
   DFF_X1 \buffer_reg[9][4][4][5]  (.D(\input_filter[4][4] [5]), .CK(n_54_15), 
      .Q(\buffer[9][4][4] [5]), .QN());
   DFF_X1 \buffer_reg[9][4][4][4]  (.D(\input_filter[4][4] [4]), .CK(n_54_15), 
      .Q(\buffer[9][4][4] [4]), .QN());
   DFF_X1 \buffer_reg[9][4][4][3]  (.D(\input_filter[4][4] [3]), .CK(n_54_15), 
      .Q(\buffer[9][4][4] [3]), .QN());
   DFF_X1 \buffer_reg[9][4][4][2]  (.D(\input_filter[4][4] [2]), .CK(n_54_15), 
      .Q(\buffer[9][4][4] [2]), .QN());
   DFF_X1 \buffer_reg[9][4][4][1]  (.D(\input_filter[4][4] [1]), .CK(n_54_15), 
      .Q(\buffer[9][4][4] [1]), .QN());
   DFF_X1 \buffer_reg[9][4][4][0]  (.D(\input_filter[4][4] [0]), .CK(n_54_15), 
      .Q(\buffer[9][4][4] [0]), .QN());
   CLKGATETST_X1 \clk_gate_buffer_reg[10][4][4]_reg  (.CK(read), .E(n_10), 
      .SE(1'b0), .GCK(n_54_0));
   DFF_X1 \buffer_reg[10][4][4][15]  (.D(\input_filter[4][4] [15]), .CK(n_54_0), 
      .Q(\buffer[10][4][4] [15]), .QN());
   DFF_X1 \buffer_reg[10][4][4][14]  (.D(\input_filter[4][4] [14]), .CK(n_54_0), 
      .Q(\buffer[10][4][4] [14]), .QN());
   DFF_X1 \buffer_reg[10][4][4][13]  (.D(\input_filter[4][4] [13]), .CK(n_54_0), 
      .Q(\buffer[10][4][4] [13]), .QN());
   DFF_X1 \buffer_reg[10][4][4][12]  (.D(\input_filter[4][4] [12]), .CK(n_54_0), 
      .Q(\buffer[10][4][4] [12]), .QN());
   DFF_X1 \buffer_reg[10][4][4][11]  (.D(\input_filter[4][4] [11]), .CK(n_54_0), 
      .Q(\buffer[10][4][4] [11]), .QN());
   DFF_X1 \buffer_reg[10][4][4][10]  (.D(\input_filter[4][4] [10]), .CK(n_54_0), 
      .Q(\buffer[10][4][4] [10]), .QN());
   DFF_X1 \buffer_reg[10][4][4][9]  (.D(\input_filter[4][4] [9]), .CK(n_54_0), 
      .Q(\buffer[10][4][4] [9]), .QN());
   DFF_X1 \buffer_reg[10][4][4][8]  (.D(\input_filter[4][4] [8]), .CK(n_54_0), 
      .Q(\buffer[10][4][4] [8]), .QN());
   DFF_X1 \buffer_reg[10][4][4][7]  (.D(\input_filter[4][4] [7]), .CK(n_54_0), 
      .Q(\buffer[10][4][4] [7]), .QN());
   DFF_X1 \buffer_reg[10][4][4][6]  (.D(\input_filter[4][4] [6]), .CK(n_54_0), 
      .Q(\buffer[10][4][4] [6]), .QN());
   DFF_X1 \buffer_reg[10][4][4][5]  (.D(\input_filter[4][4] [5]), .CK(n_54_0), 
      .Q(\buffer[10][4][4] [5]), .QN());
   DFF_X1 \buffer_reg[10][4][4][4]  (.D(\input_filter[4][4] [4]), .CK(n_54_0), 
      .Q(\buffer[10][4][4] [4]), .QN());
   DFF_X1 \buffer_reg[10][4][4][3]  (.D(\input_filter[4][4] [3]), .CK(n_54_0), 
      .Q(\buffer[10][4][4] [3]), .QN());
   DFF_X1 \buffer_reg[10][4][4][2]  (.D(\input_filter[4][4] [2]), .CK(n_54_0), 
      .Q(\buffer[10][4][4] [2]), .QN());
   DFF_X1 \buffer_reg[10][4][4][1]  (.D(\input_filter[4][4] [1]), .CK(n_54_0), 
      .Q(\buffer[10][4][4] [1]), .QN());
   DFF_X1 \buffer_reg[10][4][4][0]  (.D(\input_filter[4][4] [0]), .CK(n_54_0), 
      .Q(\buffer[10][4][4] [0]), .QN());
   CLKGATETST_X1 \clk_gate_buffer_reg[11][4][4]_reg  (.CK(read), .E(n_11), 
      .SE(1'b0), .GCK(n_54_1));
   DFF_X1 \buffer_reg[11][4][4][15]  (.D(\input_filter[4][4] [15]), .CK(n_54_1), 
      .Q(\buffer[11][4][4] [15]), .QN());
   DFF_X1 \buffer_reg[11][4][4][14]  (.D(\input_filter[4][4] [14]), .CK(n_54_1), 
      .Q(\buffer[11][4][4] [14]), .QN());
   DFF_X1 \buffer_reg[11][4][4][13]  (.D(\input_filter[4][4] [13]), .CK(n_54_1), 
      .Q(\buffer[11][4][4] [13]), .QN());
   DFF_X1 \buffer_reg[11][4][4][12]  (.D(\input_filter[4][4] [12]), .CK(n_54_1), 
      .Q(\buffer[11][4][4] [12]), .QN());
   DFF_X1 \buffer_reg[11][4][4][11]  (.D(\input_filter[4][4] [11]), .CK(n_54_1), 
      .Q(\buffer[11][4][4] [11]), .QN());
   DFF_X1 \buffer_reg[11][4][4][10]  (.D(\input_filter[4][4] [10]), .CK(n_54_1), 
      .Q(\buffer[11][4][4] [10]), .QN());
   DFF_X1 \buffer_reg[11][4][4][9]  (.D(\input_filter[4][4] [9]), .CK(n_54_1), 
      .Q(\buffer[11][4][4] [9]), .QN());
   DFF_X1 \buffer_reg[11][4][4][8]  (.D(\input_filter[4][4] [8]), .CK(n_54_1), 
      .Q(\buffer[11][4][4] [8]), .QN());
   DFF_X1 \buffer_reg[11][4][4][7]  (.D(\input_filter[4][4] [7]), .CK(n_54_1), 
      .Q(\buffer[11][4][4] [7]), .QN());
   DFF_X1 \buffer_reg[11][4][4][6]  (.D(\input_filter[4][4] [6]), .CK(n_54_1), 
      .Q(\buffer[11][4][4] [6]), .QN());
   DFF_X1 \buffer_reg[11][4][4][5]  (.D(\input_filter[4][4] [5]), .CK(n_54_1), 
      .Q(\buffer[11][4][4] [5]), .QN());
   DFF_X1 \buffer_reg[11][4][4][4]  (.D(\input_filter[4][4] [4]), .CK(n_54_1), 
      .Q(\buffer[11][4][4] [4]), .QN());
   DFF_X1 \buffer_reg[11][4][4][3]  (.D(\input_filter[4][4] [3]), .CK(n_54_1), 
      .Q(\buffer[11][4][4] [3]), .QN());
   DFF_X1 \buffer_reg[11][4][4][2]  (.D(\input_filter[4][4] [2]), .CK(n_54_1), 
      .Q(\buffer[11][4][4] [2]), .QN());
   DFF_X1 \buffer_reg[11][4][4][1]  (.D(\input_filter[4][4] [1]), .CK(n_54_1), 
      .Q(\buffer[11][4][4] [1]), .QN());
   DFF_X1 \buffer_reg[11][4][4][0]  (.D(\input_filter[4][4] [0]), .CK(n_54_1), 
      .Q(\buffer[11][4][4] [0]), .QN());
   CLKGATETST_X1 \clk_gate_buffer_reg[12][4][4]_reg  (.CK(read), .E(n_12), 
      .SE(1'b0), .GCK(n_54_2));
   DFF_X1 \buffer_reg[12][4][4][15]  (.D(\input_filter[4][4] [15]), .CK(n_54_2), 
      .Q(\buffer[12][4][4] [15]), .QN());
   DFF_X1 \buffer_reg[12][4][4][14]  (.D(\input_filter[4][4] [14]), .CK(n_54_2), 
      .Q(\buffer[12][4][4] [14]), .QN());
   DFF_X1 \buffer_reg[12][4][4][13]  (.D(\input_filter[4][4] [13]), .CK(n_54_2), 
      .Q(\buffer[12][4][4] [13]), .QN());
   DFF_X1 \buffer_reg[12][4][4][12]  (.D(\input_filter[4][4] [12]), .CK(n_54_2), 
      .Q(\buffer[12][4][4] [12]), .QN());
   DFF_X1 \buffer_reg[12][4][4][11]  (.D(\input_filter[4][4] [11]), .CK(n_54_2), 
      .Q(\buffer[12][4][4] [11]), .QN());
   DFF_X1 \buffer_reg[12][4][4][10]  (.D(\input_filter[4][4] [10]), .CK(n_54_2), 
      .Q(\buffer[12][4][4] [10]), .QN());
   DFF_X1 \buffer_reg[12][4][4][9]  (.D(\input_filter[4][4] [9]), .CK(n_54_2), 
      .Q(\buffer[12][4][4] [9]), .QN());
   DFF_X1 \buffer_reg[12][4][4][8]  (.D(\input_filter[4][4] [8]), .CK(n_54_2), 
      .Q(\buffer[12][4][4] [8]), .QN());
   DFF_X1 \buffer_reg[12][4][4][7]  (.D(\input_filter[4][4] [7]), .CK(n_54_2), 
      .Q(\buffer[12][4][4] [7]), .QN());
   DFF_X1 \buffer_reg[12][4][4][6]  (.D(\input_filter[4][4] [6]), .CK(n_54_2), 
      .Q(\buffer[12][4][4] [6]), .QN());
   DFF_X1 \buffer_reg[12][4][4][5]  (.D(\input_filter[4][4] [5]), .CK(n_54_2), 
      .Q(\buffer[12][4][4] [5]), .QN());
   DFF_X1 \buffer_reg[12][4][4][4]  (.D(\input_filter[4][4] [4]), .CK(n_54_2), 
      .Q(\buffer[12][4][4] [4]), .QN());
   DFF_X1 \buffer_reg[12][4][4][3]  (.D(\input_filter[4][4] [3]), .CK(n_54_2), 
      .Q(\buffer[12][4][4] [3]), .QN());
   DFF_X1 \buffer_reg[12][4][4][2]  (.D(\input_filter[4][4] [2]), .CK(n_54_2), 
      .Q(\buffer[12][4][4] [2]), .QN());
   DFF_X1 \buffer_reg[12][4][4][1]  (.D(\input_filter[4][4] [1]), .CK(n_54_2), 
      .Q(\buffer[12][4][4] [1]), .QN());
   DFF_X1 \buffer_reg[12][4][4][0]  (.D(\input_filter[4][4] [0]), .CK(n_54_2), 
      .Q(\buffer[12][4][4] [0]), .QN());
   DFF_X1 \buffer_reg[13][4][4][15]  (.D(\input_filter[4][4] [15]), .CK(n_54_7), 
      .Q(\buffer[13][4][4] [15]), .QN());
   DFF_X1 \buffer_reg[13][4][4][14]  (.D(\input_filter[4][4] [14]), .CK(n_54_7), 
      .Q(\buffer[13][4][4] [14]), .QN());
   DFF_X1 \buffer_reg[13][4][4][13]  (.D(\input_filter[4][4] [13]), .CK(n_54_7), 
      .Q(\buffer[13][4][4] [13]), .QN());
   DFF_X1 \buffer_reg[13][4][4][12]  (.D(\input_filter[4][4] [12]), .CK(n_54_7), 
      .Q(\buffer[13][4][4] [12]), .QN());
   DFF_X1 \buffer_reg[13][4][4][11]  (.D(\input_filter[4][4] [11]), .CK(n_54_7), 
      .Q(\buffer[13][4][4] [11]), .QN());
   DFF_X1 \buffer_reg[13][4][4][10]  (.D(\input_filter[4][4] [10]), .CK(n_54_7), 
      .Q(\buffer[13][4][4] [10]), .QN());
   DFF_X1 \buffer_reg[13][4][4][9]  (.D(\input_filter[4][4] [9]), .CK(n_54_7), 
      .Q(\buffer[13][4][4] [9]), .QN());
   DFF_X1 \buffer_reg[13][4][4][8]  (.D(\input_filter[4][4] [8]), .CK(n_54_7), 
      .Q(\buffer[13][4][4] [8]), .QN());
   DFF_X1 \buffer_reg[13][4][4][7]  (.D(\input_filter[4][4] [7]), .CK(n_54_7), 
      .Q(\buffer[13][4][4] [7]), .QN());
   DFF_X1 \buffer_reg[13][4][4][6]  (.D(\input_filter[4][4] [6]), .CK(n_54_7), 
      .Q(\buffer[13][4][4] [6]), .QN());
   DFF_X1 \buffer_reg[13][4][4][5]  (.D(\input_filter[4][4] [5]), .CK(n_54_7), 
      .Q(\buffer[13][4][4] [5]), .QN());
   DFF_X1 \buffer_reg[13][4][4][4]  (.D(\input_filter[4][4] [4]), .CK(n_54_7), 
      .Q(\buffer[13][4][4] [4]), .QN());
   DFF_X1 \buffer_reg[13][4][4][3]  (.D(\input_filter[4][4] [3]), .CK(n_54_7), 
      .Q(\buffer[13][4][4] [3]), .QN());
   DFF_X1 \buffer_reg[13][4][4][2]  (.D(\input_filter[4][4] [2]), .CK(n_54_7), 
      .Q(\buffer[13][4][4] [2]), .QN());
   DFF_X1 \buffer_reg[13][4][4][1]  (.D(\input_filter[4][4] [1]), .CK(n_54_7), 
      .Q(\buffer[13][4][4] [1]), .QN());
   DFF_X1 \buffer_reg[13][4][4][0]  (.D(\input_filter[4][4] [0]), .CK(n_54_7), 
      .Q(\buffer[13][4][4] [0]), .QN());
   DFF_X1 \buffer_reg[14][4][4][15]  (.D(\input_filter[4][4] [15]), .CK(n_54_8), 
      .Q(\buffer[14][4][4] [15]), .QN());
   DFF_X1 \buffer_reg[14][4][4][14]  (.D(\input_filter[4][4] [14]), .CK(n_54_8), 
      .Q(\buffer[14][4][4] [14]), .QN());
   DFF_X1 \buffer_reg[14][4][4][13]  (.D(\input_filter[4][4] [13]), .CK(n_54_8), 
      .Q(\buffer[14][4][4] [13]), .QN());
   DFF_X1 \buffer_reg[14][4][4][12]  (.D(\input_filter[4][4] [12]), .CK(n_54_8), 
      .Q(\buffer[14][4][4] [12]), .QN());
   DFF_X1 \buffer_reg[14][4][4][11]  (.D(\input_filter[4][4] [11]), .CK(n_54_8), 
      .Q(\buffer[14][4][4] [11]), .QN());
   DFF_X1 \buffer_reg[14][4][4][10]  (.D(\input_filter[4][4] [10]), .CK(n_54_8), 
      .Q(\buffer[14][4][4] [10]), .QN());
   DFF_X1 \buffer_reg[14][4][4][9]  (.D(\input_filter[4][4] [9]), .CK(n_54_8), 
      .Q(\buffer[14][4][4] [9]), .QN());
   DFF_X1 \buffer_reg[14][4][4][8]  (.D(\input_filter[4][4] [8]), .CK(n_54_8), 
      .Q(\buffer[14][4][4] [8]), .QN());
   DFF_X1 \buffer_reg[14][4][4][7]  (.D(\input_filter[4][4] [7]), .CK(n_54_8), 
      .Q(\buffer[14][4][4] [7]), .QN());
   DFF_X1 \buffer_reg[14][4][4][6]  (.D(\input_filter[4][4] [6]), .CK(n_54_8), 
      .Q(\buffer[14][4][4] [6]), .QN());
   DFF_X1 \buffer_reg[14][4][4][5]  (.D(\input_filter[4][4] [5]), .CK(n_54_8), 
      .Q(\buffer[14][4][4] [5]), .QN());
   DFF_X1 \buffer_reg[14][4][4][4]  (.D(\input_filter[4][4] [4]), .CK(n_54_8), 
      .Q(\buffer[14][4][4] [4]), .QN());
   DFF_X1 \buffer_reg[14][4][4][3]  (.D(\input_filter[4][4] [3]), .CK(n_54_8), 
      .Q(\buffer[14][4][4] [3]), .QN());
   DFF_X1 \buffer_reg[14][4][4][2]  (.D(\input_filter[4][4] [2]), .CK(n_54_8), 
      .Q(\buffer[14][4][4] [2]), .QN());
   DFF_X1 \buffer_reg[14][4][4][1]  (.D(\input_filter[4][4] [1]), .CK(n_54_8), 
      .Q(\buffer[14][4][4] [1]), .QN());
   DFF_X1 \buffer_reg[14][4][4][0]  (.D(\input_filter[4][4] [0]), .CK(n_54_8), 
      .Q(\buffer[14][4][4] [0]), .QN());
   DFF_X1 \buffer_reg[15][4][4][15]  (.D(\input_filter[4][4] [15]), .CK(n_54_9), 
      .Q(\buffer[15][4][4] [15]), .QN());
   DFF_X1 \buffer_reg[15][4][4][14]  (.D(\input_filter[4][4] [14]), .CK(n_54_9), 
      .Q(\buffer[15][4][4] [14]), .QN());
   DFF_X1 \buffer_reg[15][4][4][13]  (.D(\input_filter[4][4] [13]), .CK(n_54_9), 
      .Q(\buffer[15][4][4] [13]), .QN());
   DFF_X1 \buffer_reg[15][4][4][12]  (.D(\input_filter[4][4] [12]), .CK(n_54_9), 
      .Q(\buffer[15][4][4] [12]), .QN());
   DFF_X1 \buffer_reg[15][4][4][11]  (.D(\input_filter[4][4] [11]), .CK(n_54_9), 
      .Q(\buffer[15][4][4] [11]), .QN());
   DFF_X1 \buffer_reg[15][4][4][10]  (.D(\input_filter[4][4] [10]), .CK(n_54_9), 
      .Q(\buffer[15][4][4] [10]), .QN());
   DFF_X1 \buffer_reg[15][4][4][9]  (.D(\input_filter[4][4] [9]), .CK(n_54_9), 
      .Q(\buffer[15][4][4] [9]), .QN());
   DFF_X1 \buffer_reg[15][4][4][8]  (.D(\input_filter[4][4] [8]), .CK(n_54_9), 
      .Q(\buffer[15][4][4] [8]), .QN());
   DFF_X1 \buffer_reg[15][4][4][7]  (.D(\input_filter[4][4] [7]), .CK(n_54_9), 
      .Q(\buffer[15][4][4] [7]), .QN());
   DFF_X1 \buffer_reg[15][4][4][6]  (.D(\input_filter[4][4] [6]), .CK(n_54_9), 
      .Q(\buffer[15][4][4] [6]), .QN());
   DFF_X1 \buffer_reg[15][4][4][5]  (.D(\input_filter[4][4] [5]), .CK(n_54_9), 
      .Q(\buffer[15][4][4] [5]), .QN());
   DFF_X1 \buffer_reg[15][4][4][4]  (.D(\input_filter[4][4] [4]), .CK(n_54_9), 
      .Q(\buffer[15][4][4] [4]), .QN());
   DFF_X1 \buffer_reg[15][4][4][3]  (.D(\input_filter[4][4] [3]), .CK(n_54_9), 
      .Q(\buffer[15][4][4] [3]), .QN());
   DFF_X1 \buffer_reg[15][4][4][2]  (.D(\input_filter[4][4] [2]), .CK(n_54_9), 
      .Q(\buffer[15][4][4] [2]), .QN());
   DFF_X1 \buffer_reg[15][4][4][1]  (.D(\input_filter[4][4] [1]), .CK(n_54_9), 
      .Q(\buffer[15][4][4] [1]), .QN());
   DFF_X1 \buffer_reg[15][4][4][0]  (.D(\input_filter[4][4] [0]), .CK(n_54_9), 
      .Q(\buffer[15][4][4] [0]), .QN());
   DFF_X1 \buffer_reg[15][0][0][15]  (.D(\input_filter[0][0] [15]), .CK(n_54_9), 
      .Q(\buffer[15][0][0] [15]), .QN());
   DFF_X1 \buffer_reg[15][0][0][14]  (.D(\input_filter[0][0] [14]), .CK(n_54_9), 
      .Q(\buffer[15][0][0] [14]), .QN());
   DFF_X1 \buffer_reg[15][0][0][13]  (.D(\input_filter[0][0] [13]), .CK(n_54_9), 
      .Q(\buffer[15][0][0] [13]), .QN());
   DFF_X1 \buffer_reg[15][0][0][12]  (.D(\input_filter[0][0] [12]), .CK(n_54_9), 
      .Q(\buffer[15][0][0] [12]), .QN());
   DFF_X1 \buffer_reg[15][0][0][11]  (.D(\input_filter[0][0] [11]), .CK(n_54_9), 
      .Q(\buffer[15][0][0] [11]), .QN());
   DFF_X1 \buffer_reg[15][0][0][10]  (.D(\input_filter[0][0] [10]), .CK(n_54_9), 
      .Q(\buffer[15][0][0] [10]), .QN());
   DFF_X1 \buffer_reg[15][0][0][9]  (.D(\input_filter[0][0] [9]), .CK(n_54_9), 
      .Q(\buffer[15][0][0] [9]), .QN());
   DFF_X1 \buffer_reg[15][0][0][8]  (.D(\input_filter[0][0] [8]), .CK(n_54_9), 
      .Q(\buffer[15][0][0] [8]), .QN());
   DFF_X1 \buffer_reg[15][0][0][7]  (.D(\input_filter[0][0] [7]), .CK(n_54_9), 
      .Q(\buffer[15][0][0] [7]), .QN());
   DFF_X1 \buffer_reg[15][0][0][6]  (.D(\input_filter[0][0] [6]), .CK(n_54_9), 
      .Q(\buffer[15][0][0] [6]), .QN());
   DFF_X1 \buffer_reg[15][0][0][5]  (.D(\input_filter[0][0] [5]), .CK(n_54_9), 
      .Q(\buffer[15][0][0] [5]), .QN());
   DFF_X1 \buffer_reg[15][0][0][4]  (.D(\input_filter[0][0] [4]), .CK(n_54_9), 
      .Q(\buffer[15][0][0] [4]), .QN());
   DFF_X1 \buffer_reg[15][0][0][3]  (.D(\input_filter[0][0] [3]), .CK(n_54_9), 
      .Q(\buffer[15][0][0] [3]), .QN());
   DFF_X1 \buffer_reg[15][0][0][2]  (.D(\input_filter[0][0] [2]), .CK(n_54_9), 
      .Q(\buffer[15][0][0] [2]), .QN());
   DFF_X1 \buffer_reg[15][0][0][1]  (.D(\input_filter[0][0] [1]), .CK(n_54_9), 
      .Q(\buffer[15][0][0] [1]), .QN());
   DFF_X1 \buffer_reg[15][0][0][0]  (.D(\input_filter[0][0] [0]), .CK(n_54_9), 
      .Q(\buffer[15][0][0] [0]), .QN());
   DFF_X1 \buffer_reg[2][0][0][15]  (.D(\input_filter[0][0] [15]), .CK(n_54_4), 
      .Q(\buffer[2][0][0] [15]), .QN());
   DFF_X1 \buffer_reg[2][0][0][14]  (.D(\input_filter[0][0] [14]), .CK(n_54_4), 
      .Q(\buffer[2][0][0] [14]), .QN());
   DFF_X1 \buffer_reg[2][0][0][13]  (.D(\input_filter[0][0] [13]), .CK(n_54_4), 
      .Q(\buffer[2][0][0] [13]), .QN());
   DFF_X1 \buffer_reg[2][0][0][12]  (.D(\input_filter[0][0] [12]), .CK(n_54_4), 
      .Q(\buffer[2][0][0] [12]), .QN());
   DFF_X1 \buffer_reg[2][0][0][11]  (.D(\input_filter[0][0] [11]), .CK(n_54_4), 
      .Q(\buffer[2][0][0] [11]), .QN());
   DFF_X1 \buffer_reg[2][0][0][10]  (.D(\input_filter[0][0] [10]), .CK(n_54_4), 
      .Q(\buffer[2][0][0] [10]), .QN());
   DFF_X1 \buffer_reg[2][0][0][9]  (.D(\input_filter[0][0] [9]), .CK(n_54_4), 
      .Q(\buffer[2][0][0] [9]), .QN());
   DFF_X1 \buffer_reg[2][0][0][8]  (.D(\input_filter[0][0] [8]), .CK(n_54_4), 
      .Q(\buffer[2][0][0] [8]), .QN());
   DFF_X1 \buffer_reg[2][0][0][7]  (.D(\input_filter[0][0] [7]), .CK(n_54_4), 
      .Q(\buffer[2][0][0] [7]), .QN());
   DFF_X1 \buffer_reg[2][0][0][6]  (.D(\input_filter[0][0] [6]), .CK(n_54_4), 
      .Q(\buffer[2][0][0] [6]), .QN());
   DFF_X1 \buffer_reg[2][0][0][5]  (.D(\input_filter[0][0] [5]), .CK(n_54_4), 
      .Q(\buffer[2][0][0] [5]), .QN());
   DFF_X1 \buffer_reg[2][0][0][4]  (.D(\input_filter[0][0] [4]), .CK(n_54_4), 
      .Q(\buffer[2][0][0] [4]), .QN());
   DFF_X1 \buffer_reg[2][0][0][3]  (.D(\input_filter[0][0] [3]), .CK(n_54_4), 
      .Q(\buffer[2][0][0] [3]), .QN());
   DFF_X1 \buffer_reg[2][0][0][2]  (.D(\input_filter[0][0] [2]), .CK(n_54_4), 
      .Q(\buffer[2][0][0] [2]), .QN());
   DFF_X1 \buffer_reg[2][0][0][1]  (.D(\input_filter[0][0] [1]), .CK(n_54_4), 
      .Q(\buffer[2][0][0] [1]), .QN());
   DFF_X1 \buffer_reg[2][0][0][0]  (.D(\input_filter[0][0] [0]), .CK(n_54_4), 
      .Q(\buffer[2][0][0] [0]), .QN());
   DFF_X1 \buffer_reg[1][0][0][15]  (.D(\input_filter[0][0] [15]), .CK(n_54_3), 
      .Q(\buffer[1][0][0] [15]), .QN());
   DFF_X1 \buffer_reg[1][0][0][14]  (.D(\input_filter[0][0] [14]), .CK(n_54_3), 
      .Q(\buffer[1][0][0] [14]), .QN());
   DFF_X1 \buffer_reg[1][0][0][13]  (.D(\input_filter[0][0] [13]), .CK(n_54_3), 
      .Q(\buffer[1][0][0] [13]), .QN());
   DFF_X1 \buffer_reg[1][0][0][12]  (.D(\input_filter[0][0] [12]), .CK(n_54_3), 
      .Q(\buffer[1][0][0] [12]), .QN());
   DFF_X1 \buffer_reg[1][0][0][11]  (.D(\input_filter[0][0] [11]), .CK(n_54_3), 
      .Q(\buffer[1][0][0] [11]), .QN());
   DFF_X1 \buffer_reg[1][0][0][10]  (.D(\input_filter[0][0] [10]), .CK(n_54_3), 
      .Q(\buffer[1][0][0] [10]), .QN());
   DFF_X1 \buffer_reg[1][0][0][9]  (.D(\input_filter[0][0] [9]), .CK(n_54_3), 
      .Q(\buffer[1][0][0] [9]), .QN());
   DFF_X1 \buffer_reg[1][0][0][8]  (.D(\input_filter[0][0] [8]), .CK(n_54_3), 
      .Q(\buffer[1][0][0] [8]), .QN());
   DFF_X1 \buffer_reg[1][0][0][7]  (.D(\input_filter[0][0] [7]), .CK(n_54_3), 
      .Q(\buffer[1][0][0] [7]), .QN());
   DFF_X1 \buffer_reg[1][0][0][6]  (.D(\input_filter[0][0] [6]), .CK(n_54_3), 
      .Q(\buffer[1][0][0] [6]), .QN());
   DFF_X1 \buffer_reg[1][0][0][5]  (.D(\input_filter[0][0] [5]), .CK(n_54_3), 
      .Q(\buffer[1][0][0] [5]), .QN());
   DFF_X1 \buffer_reg[1][0][0][4]  (.D(\input_filter[0][0] [4]), .CK(n_54_3), 
      .Q(\buffer[1][0][0] [4]), .QN());
   DFF_X1 \buffer_reg[1][0][0][3]  (.D(\input_filter[0][0] [3]), .CK(n_54_3), 
      .Q(\buffer[1][0][0] [3]), .QN());
   DFF_X1 \buffer_reg[1][0][0][2]  (.D(\input_filter[0][0] [2]), .CK(n_54_3), 
      .Q(\buffer[1][0][0] [2]), .QN());
   DFF_X1 \buffer_reg[1][0][0][1]  (.D(\input_filter[0][0] [1]), .CK(n_54_3), 
      .Q(\buffer[1][0][0] [1]), .QN());
   DFF_X1 \buffer_reg[1][0][0][0]  (.D(\input_filter[0][0] [0]), .CK(n_54_3), 
      .Q(\buffer[1][0][0] [0]), .QN());
   CLKGATETST_X1 \clk_gate_buffer_reg[1][4][3]_reg  (.CK(read), .E(n_1), 
      .SE(1'b0), .GCK(n_54_3));
   CLKGATETST_X1 \clk_gate_buffer_reg[2][4][3]_reg  (.CK(read), .E(n_2), 
      .SE(1'b0), .GCK(n_54_4));
   CLKGATETST_X1 \clk_gate_buffer_reg[3][4][3]_reg  (.CK(read), .E(n_3), 
      .SE(1'b0), .GCK(n_54_5));
   CLKGATETST_X1 \clk_gate_buffer_reg[13][4][3]_reg  (.CK(read), .E(n_13), 
      .SE(1'b0), .GCK(n_54_7));
   CLKGATETST_X1 \clk_gate_buffer_reg[14][4][3]_reg  (.CK(read), .E(n_14), 
      .SE(1'b0), .GCK(n_54_8));
   CLKGATETST_X1 \clk_gate_buffer_reg[15][4][3]_reg  (.CK(read), .E(n_15), 
      .SE(1'b0), .GCK(n_54_9));
   DFF_X1 \buffer_reg[12][3][2][15]  (.D(\input_filter[3][2] [15]), .CK(n_55_0), 
      .Q(\buffer[12][3][2] [15]), .QN());
   DFF_X1 \buffer_reg[12][3][2][14]  (.D(\input_filter[3][2] [14]), .CK(n_55_0), 
      .Q(\buffer[12][3][2] [14]), .QN());
   DFF_X1 \buffer_reg[12][3][2][13]  (.D(\input_filter[3][2] [13]), .CK(n_55_0), 
      .Q(\buffer[12][3][2] [13]), .QN());
   DFF_X1 \buffer_reg[12][3][2][12]  (.D(\input_filter[3][2] [12]), .CK(n_55_0), 
      .Q(\buffer[12][3][2] [12]), .QN());
   DFF_X1 \buffer_reg[12][3][2][11]  (.D(\input_filter[3][2] [11]), .CK(n_55_0), 
      .Q(\buffer[12][3][2] [11]), .QN());
   DFF_X1 \buffer_reg[12][3][2][10]  (.D(\input_filter[3][2] [10]), .CK(n_55_0), 
      .Q(\buffer[12][3][2] [10]), .QN());
   DFF_X1 \buffer_reg[12][3][2][9]  (.D(\input_filter[3][2] [9]), .CK(n_55_0), 
      .Q(\buffer[12][3][2] [9]), .QN());
   DFF_X1 \buffer_reg[12][3][2][8]  (.D(\input_filter[3][2] [8]), .CK(n_55_0), 
      .Q(\buffer[12][3][2] [8]), .QN());
   DFF_X1 \buffer_reg[12][3][2][7]  (.D(\input_filter[3][2] [7]), .CK(n_55_0), 
      .Q(\buffer[12][3][2] [7]), .QN());
   DFF_X1 \buffer_reg[12][3][2][6]  (.D(\input_filter[3][2] [6]), .CK(n_55_0), 
      .Q(\buffer[12][3][2] [6]), .QN());
   DFF_X1 \buffer_reg[12][3][2][5]  (.D(\input_filter[3][2] [5]), .CK(n_55_0), 
      .Q(\buffer[12][3][2] [5]), .QN());
   DFF_X1 \buffer_reg[12][3][2][4]  (.D(\input_filter[3][2] [4]), .CK(n_55_0), 
      .Q(\buffer[12][3][2] [4]), .QN());
   DFF_X1 \buffer_reg[12][3][2][3]  (.D(\input_filter[3][2] [3]), .CK(n_55_0), 
      .Q(\buffer[12][3][2] [3]), .QN());
   DFF_X1 \buffer_reg[12][3][2][2]  (.D(\input_filter[3][2] [2]), .CK(n_55_0), 
      .Q(\buffer[12][3][2] [2]), .QN());
   DFF_X1 \buffer_reg[12][3][2][1]  (.D(\input_filter[3][2] [1]), .CK(n_55_0), 
      .Q(\buffer[12][3][2] [1]), .QN());
   DFF_X1 \buffer_reg[12][3][2][0]  (.D(\input_filter[3][2] [0]), .CK(n_55_0), 
      .Q(\buffer[12][3][2] [0]), .QN());
   DFF_X1 \buffer_reg[11][3][2][15]  (.D(\input_filter[3][2] [15]), .CK(n_55_1), 
      .Q(\buffer[11][3][2] [15]), .QN());
   DFF_X1 \buffer_reg[11][3][2][14]  (.D(\input_filter[3][2] [14]), .CK(n_55_1), 
      .Q(\buffer[11][3][2] [14]), .QN());
   DFF_X1 \buffer_reg[11][3][2][13]  (.D(\input_filter[3][2] [13]), .CK(n_55_1), 
      .Q(\buffer[11][3][2] [13]), .QN());
   DFF_X1 \buffer_reg[11][3][2][12]  (.D(\input_filter[3][2] [12]), .CK(n_55_1), 
      .Q(\buffer[11][3][2] [12]), .QN());
   DFF_X1 \buffer_reg[11][3][2][11]  (.D(\input_filter[3][2] [11]), .CK(n_55_1), 
      .Q(\buffer[11][3][2] [11]), .QN());
   DFF_X1 \buffer_reg[11][3][2][10]  (.D(\input_filter[3][2] [10]), .CK(n_55_1), 
      .Q(\buffer[11][3][2] [10]), .QN());
   DFF_X1 \buffer_reg[11][3][2][9]  (.D(\input_filter[3][2] [9]), .CK(n_55_1), 
      .Q(\buffer[11][3][2] [9]), .QN());
   DFF_X1 \buffer_reg[11][3][2][8]  (.D(\input_filter[3][2] [8]), .CK(n_55_1), 
      .Q(\buffer[11][3][2] [8]), .QN());
   DFF_X1 \buffer_reg[11][3][2][7]  (.D(\input_filter[3][2] [7]), .CK(n_55_1), 
      .Q(\buffer[11][3][2] [7]), .QN());
   DFF_X1 \buffer_reg[11][3][2][6]  (.D(\input_filter[3][2] [6]), .CK(n_55_1), 
      .Q(\buffer[11][3][2] [6]), .QN());
   DFF_X1 \buffer_reg[11][3][2][5]  (.D(\input_filter[3][2] [5]), .CK(n_55_1), 
      .Q(\buffer[11][3][2] [5]), .QN());
   DFF_X1 \buffer_reg[11][3][2][4]  (.D(\input_filter[3][2] [4]), .CK(n_55_1), 
      .Q(\buffer[11][3][2] [4]), .QN());
   DFF_X1 \buffer_reg[11][3][2][3]  (.D(\input_filter[3][2] [3]), .CK(n_55_1), 
      .Q(\buffer[11][3][2] [3]), .QN());
   DFF_X1 \buffer_reg[11][3][2][2]  (.D(\input_filter[3][2] [2]), .CK(n_55_1), 
      .Q(\buffer[11][3][2] [2]), .QN());
   DFF_X1 \buffer_reg[11][3][2][1]  (.D(\input_filter[3][2] [1]), .CK(n_55_1), 
      .Q(\buffer[11][3][2] [1]), .QN());
   DFF_X1 \buffer_reg[11][3][2][0]  (.D(\input_filter[3][2] [0]), .CK(n_55_1), 
      .Q(\buffer[11][3][2] [0]), .QN());
   DFF_X1 \buffer_reg[10][3][2][15]  (.D(\input_filter[3][2] [15]), .CK(n_55_2), 
      .Q(\buffer[10][3][2] [15]), .QN());
   DFF_X1 \buffer_reg[10][3][2][14]  (.D(\input_filter[3][2] [14]), .CK(n_55_2), 
      .Q(\buffer[10][3][2] [14]), .QN());
   DFF_X1 \buffer_reg[10][3][2][13]  (.D(\input_filter[3][2] [13]), .CK(n_55_2), 
      .Q(\buffer[10][3][2] [13]), .QN());
   DFF_X1 \buffer_reg[10][3][2][12]  (.D(\input_filter[3][2] [12]), .CK(n_55_2), 
      .Q(\buffer[10][3][2] [12]), .QN());
   DFF_X1 \buffer_reg[10][3][2][11]  (.D(\input_filter[3][2] [11]), .CK(n_55_2), 
      .Q(\buffer[10][3][2] [11]), .QN());
   DFF_X1 \buffer_reg[10][3][2][10]  (.D(\input_filter[3][2] [10]), .CK(n_55_2), 
      .Q(\buffer[10][3][2] [10]), .QN());
   DFF_X1 \buffer_reg[10][3][2][9]  (.D(\input_filter[3][2] [9]), .CK(n_55_2), 
      .Q(\buffer[10][3][2] [9]), .QN());
   DFF_X1 \buffer_reg[10][3][2][8]  (.D(\input_filter[3][2] [8]), .CK(n_55_2), 
      .Q(\buffer[10][3][2] [8]), .QN());
   DFF_X1 \buffer_reg[10][3][2][7]  (.D(\input_filter[3][2] [7]), .CK(n_55_2), 
      .Q(\buffer[10][3][2] [7]), .QN());
   DFF_X1 \buffer_reg[10][3][2][6]  (.D(\input_filter[3][2] [6]), .CK(n_55_2), 
      .Q(\buffer[10][3][2] [6]), .QN());
   DFF_X1 \buffer_reg[10][3][2][5]  (.D(\input_filter[3][2] [5]), .CK(n_55_2), 
      .Q(\buffer[10][3][2] [5]), .QN());
   DFF_X1 \buffer_reg[10][3][2][4]  (.D(\input_filter[3][2] [4]), .CK(n_55_2), 
      .Q(\buffer[10][3][2] [4]), .QN());
   DFF_X1 \buffer_reg[10][3][2][3]  (.D(\input_filter[3][2] [3]), .CK(n_55_2), 
      .Q(\buffer[10][3][2] [3]), .QN());
   DFF_X1 \buffer_reg[10][3][2][2]  (.D(\input_filter[3][2] [2]), .CK(n_55_2), 
      .Q(\buffer[10][3][2] [2]), .QN());
   DFF_X1 \buffer_reg[10][3][2][1]  (.D(\input_filter[3][2] [1]), .CK(n_55_2), 
      .Q(\buffer[10][3][2] [1]), .QN());
   DFF_X1 \buffer_reg[10][3][2][0]  (.D(\input_filter[3][2] [0]), .CK(n_55_2), 
      .Q(\buffer[10][3][2] [0]), .QN());
   DFF_X1 \buffer_reg[9][3][2][15]  (.D(\input_filter[3][2] [15]), .CK(n_55_3), 
      .Q(\buffer[9][3][2] [15]), .QN());
   DFF_X1 \buffer_reg[9][3][2][14]  (.D(\input_filter[3][2] [14]), .CK(n_55_3), 
      .Q(\buffer[9][3][2] [14]), .QN());
   DFF_X1 \buffer_reg[9][3][2][13]  (.D(\input_filter[3][2] [13]), .CK(n_55_3), 
      .Q(\buffer[9][3][2] [13]), .QN());
   DFF_X1 \buffer_reg[9][3][2][12]  (.D(\input_filter[3][2] [12]), .CK(n_55_3), 
      .Q(\buffer[9][3][2] [12]), .QN());
   DFF_X1 \buffer_reg[9][3][2][11]  (.D(\input_filter[3][2] [11]), .CK(n_55_3), 
      .Q(\buffer[9][3][2] [11]), .QN());
   DFF_X1 \buffer_reg[9][3][2][10]  (.D(\input_filter[3][2] [10]), .CK(n_55_3), 
      .Q(\buffer[9][3][2] [10]), .QN());
   DFF_X1 \buffer_reg[9][3][2][9]  (.D(\input_filter[3][2] [9]), .CK(n_55_3), 
      .Q(\buffer[9][3][2] [9]), .QN());
   DFF_X1 \buffer_reg[9][3][2][8]  (.D(\input_filter[3][2] [8]), .CK(n_55_3), 
      .Q(\buffer[9][3][2] [8]), .QN());
   DFF_X1 \buffer_reg[9][3][2][7]  (.D(\input_filter[3][2] [7]), .CK(n_55_3), 
      .Q(\buffer[9][3][2] [7]), .QN());
   DFF_X1 \buffer_reg[9][3][2][6]  (.D(\input_filter[3][2] [6]), .CK(n_55_3), 
      .Q(\buffer[9][3][2] [6]), .QN());
   DFF_X1 \buffer_reg[9][3][2][5]  (.D(\input_filter[3][2] [5]), .CK(n_55_3), 
      .Q(\buffer[9][3][2] [5]), .QN());
   DFF_X1 \buffer_reg[9][3][2][4]  (.D(\input_filter[3][2] [4]), .CK(n_55_3), 
      .Q(\buffer[9][3][2] [4]), .QN());
   DFF_X1 \buffer_reg[9][3][2][3]  (.D(\input_filter[3][2] [3]), .CK(n_55_3), 
      .Q(\buffer[9][3][2] [3]), .QN());
   DFF_X1 \buffer_reg[9][3][2][2]  (.D(\input_filter[3][2] [2]), .CK(n_55_3), 
      .Q(\buffer[9][3][2] [2]), .QN());
   DFF_X1 \buffer_reg[9][3][2][1]  (.D(\input_filter[3][2] [1]), .CK(n_55_3), 
      .Q(\buffer[9][3][2] [1]), .QN());
   DFF_X1 \buffer_reg[9][3][2][0]  (.D(\input_filter[3][2] [0]), .CK(n_55_3), 
      .Q(\buffer[9][3][2] [0]), .QN());
   DFF_X1 \buffer_reg[8][3][2][15]  (.D(\input_filter[3][2] [15]), .CK(n_55_4), 
      .Q(\buffer[8][3][2] [15]), .QN());
   DFF_X1 \buffer_reg[8][3][2][14]  (.D(\input_filter[3][2] [14]), .CK(n_55_4), 
      .Q(\buffer[8][3][2] [14]), .QN());
   DFF_X1 \buffer_reg[8][3][2][13]  (.D(\input_filter[3][2] [13]), .CK(n_55_4), 
      .Q(\buffer[8][3][2] [13]), .QN());
   DFF_X1 \buffer_reg[8][3][2][12]  (.D(\input_filter[3][2] [12]), .CK(n_55_4), 
      .Q(\buffer[8][3][2] [12]), .QN());
   DFF_X1 \buffer_reg[8][3][2][11]  (.D(\input_filter[3][2] [11]), .CK(n_55_4), 
      .Q(\buffer[8][3][2] [11]), .QN());
   DFF_X1 \buffer_reg[8][3][2][10]  (.D(\input_filter[3][2] [10]), .CK(n_55_4), 
      .Q(\buffer[8][3][2] [10]), .QN());
   DFF_X1 \buffer_reg[8][3][2][9]  (.D(\input_filter[3][2] [9]), .CK(n_55_4), 
      .Q(\buffer[8][3][2] [9]), .QN());
   DFF_X1 \buffer_reg[8][3][2][8]  (.D(\input_filter[3][2] [8]), .CK(n_55_4), 
      .Q(\buffer[8][3][2] [8]), .QN());
   DFF_X1 \buffer_reg[8][3][2][7]  (.D(\input_filter[3][2] [7]), .CK(n_55_4), 
      .Q(\buffer[8][3][2] [7]), .QN());
   DFF_X1 \buffer_reg[8][3][2][6]  (.D(\input_filter[3][2] [6]), .CK(n_55_4), 
      .Q(\buffer[8][3][2] [6]), .QN());
   DFF_X1 \buffer_reg[8][3][2][5]  (.D(\input_filter[3][2] [5]), .CK(n_55_4), 
      .Q(\buffer[8][3][2] [5]), .QN());
   DFF_X1 \buffer_reg[8][3][2][4]  (.D(\input_filter[3][2] [4]), .CK(n_55_4), 
      .Q(\buffer[8][3][2] [4]), .QN());
   DFF_X1 \buffer_reg[8][3][2][3]  (.D(\input_filter[3][2] [3]), .CK(n_55_4), 
      .Q(\buffer[8][3][2] [3]), .QN());
   DFF_X1 \buffer_reg[8][3][2][2]  (.D(\input_filter[3][2] [2]), .CK(n_55_4), 
      .Q(\buffer[8][3][2] [2]), .QN());
   DFF_X1 \buffer_reg[8][3][2][1]  (.D(\input_filter[3][2] [1]), .CK(n_55_4), 
      .Q(\buffer[8][3][2] [1]), .QN());
   DFF_X1 \buffer_reg[8][3][2][0]  (.D(\input_filter[3][2] [0]), .CK(n_55_4), 
      .Q(\buffer[8][3][2] [0]), .QN());
   DFF_X1 \buffer_reg[7][3][2][15]  (.D(\input_filter[3][2] [15]), .CK(n_55_5), 
      .Q(\buffer[7][3][2] [15]), .QN());
   DFF_X1 \buffer_reg[7][3][2][14]  (.D(\input_filter[3][2] [14]), .CK(n_55_5), 
      .Q(\buffer[7][3][2] [14]), .QN());
   DFF_X1 \buffer_reg[7][3][2][13]  (.D(\input_filter[3][2] [13]), .CK(n_55_5), 
      .Q(\buffer[7][3][2] [13]), .QN());
   DFF_X1 \buffer_reg[7][3][2][12]  (.D(\input_filter[3][2] [12]), .CK(n_55_5), 
      .Q(\buffer[7][3][2] [12]), .QN());
   DFF_X1 \buffer_reg[7][3][2][11]  (.D(\input_filter[3][2] [11]), .CK(n_55_5), 
      .Q(\buffer[7][3][2] [11]), .QN());
   DFF_X1 \buffer_reg[7][3][2][10]  (.D(\input_filter[3][2] [10]), .CK(n_55_5), 
      .Q(\buffer[7][3][2] [10]), .QN());
   DFF_X1 \buffer_reg[7][3][2][9]  (.D(\input_filter[3][2] [9]), .CK(n_55_5), 
      .Q(\buffer[7][3][2] [9]), .QN());
   DFF_X1 \buffer_reg[7][3][2][8]  (.D(\input_filter[3][2] [8]), .CK(n_55_5), 
      .Q(\buffer[7][3][2] [8]), .QN());
   DFF_X1 \buffer_reg[7][3][2][7]  (.D(\input_filter[3][2] [7]), .CK(n_55_5), 
      .Q(\buffer[7][3][2] [7]), .QN());
   DFF_X1 \buffer_reg[7][3][2][6]  (.D(\input_filter[3][2] [6]), .CK(n_55_5), 
      .Q(\buffer[7][3][2] [6]), .QN());
   DFF_X1 \buffer_reg[7][3][2][5]  (.D(\input_filter[3][2] [5]), .CK(n_55_5), 
      .Q(\buffer[7][3][2] [5]), .QN());
   DFF_X1 \buffer_reg[7][3][2][4]  (.D(\input_filter[3][2] [4]), .CK(n_55_5), 
      .Q(\buffer[7][3][2] [4]), .QN());
   DFF_X1 \buffer_reg[7][3][2][3]  (.D(\input_filter[3][2] [3]), .CK(n_55_5), 
      .Q(\buffer[7][3][2] [3]), .QN());
   DFF_X1 \buffer_reg[7][3][2][2]  (.D(\input_filter[3][2] [2]), .CK(n_55_5), 
      .Q(\buffer[7][3][2] [2]), .QN());
   DFF_X1 \buffer_reg[7][3][2][1]  (.D(\input_filter[3][2] [1]), .CK(n_55_5), 
      .Q(\buffer[7][3][2] [1]), .QN());
   DFF_X1 \buffer_reg[7][3][2][0]  (.D(\input_filter[3][2] [0]), .CK(n_55_5), 
      .Q(\buffer[7][3][2] [0]), .QN());
   DFF_X1 \buffer_reg[6][3][2][15]  (.D(\input_filter[3][2] [15]), .CK(n_55_6), 
      .Q(\buffer[6][3][2] [15]), .QN());
   DFF_X1 \buffer_reg[6][3][2][14]  (.D(\input_filter[3][2] [14]), .CK(n_55_6), 
      .Q(\buffer[6][3][2] [14]), .QN());
   DFF_X1 \buffer_reg[6][3][2][13]  (.D(\input_filter[3][2] [13]), .CK(n_55_6), 
      .Q(\buffer[6][3][2] [13]), .QN());
   DFF_X1 \buffer_reg[6][3][2][12]  (.D(\input_filter[3][2] [12]), .CK(n_55_6), 
      .Q(\buffer[6][3][2] [12]), .QN());
   DFF_X1 \buffer_reg[6][3][2][11]  (.D(\input_filter[3][2] [11]), .CK(n_55_6), 
      .Q(\buffer[6][3][2] [11]), .QN());
   DFF_X1 \buffer_reg[6][3][2][10]  (.D(\input_filter[3][2] [10]), .CK(n_55_6), 
      .Q(\buffer[6][3][2] [10]), .QN());
   DFF_X1 \buffer_reg[6][3][2][9]  (.D(\input_filter[3][2] [9]), .CK(n_55_6), 
      .Q(\buffer[6][3][2] [9]), .QN());
   DFF_X1 \buffer_reg[6][3][2][8]  (.D(\input_filter[3][2] [8]), .CK(n_55_6), 
      .Q(\buffer[6][3][2] [8]), .QN());
   DFF_X1 \buffer_reg[6][3][2][7]  (.D(\input_filter[3][2] [7]), .CK(n_55_6), 
      .Q(\buffer[6][3][2] [7]), .QN());
   DFF_X1 \buffer_reg[6][3][2][6]  (.D(\input_filter[3][2] [6]), .CK(n_55_6), 
      .Q(\buffer[6][3][2] [6]), .QN());
   DFF_X1 \buffer_reg[6][3][2][5]  (.D(\input_filter[3][2] [5]), .CK(n_55_6), 
      .Q(\buffer[6][3][2] [5]), .QN());
   DFF_X1 \buffer_reg[6][3][2][4]  (.D(\input_filter[3][2] [4]), .CK(n_55_6), 
      .Q(\buffer[6][3][2] [4]), .QN());
   DFF_X1 \buffer_reg[6][3][2][3]  (.D(\input_filter[3][2] [3]), .CK(n_55_6), 
      .Q(\buffer[6][3][2] [3]), .QN());
   DFF_X1 \buffer_reg[6][3][2][2]  (.D(\input_filter[3][2] [2]), .CK(n_55_6), 
      .Q(\buffer[6][3][2] [2]), .QN());
   DFF_X1 \buffer_reg[6][3][2][1]  (.D(\input_filter[3][2] [1]), .CK(n_55_6), 
      .Q(\buffer[6][3][2] [1]), .QN());
   DFF_X1 \buffer_reg[6][3][2][0]  (.D(\input_filter[3][2] [0]), .CK(n_55_6), 
      .Q(\buffer[6][3][2] [0]), .QN());
   DFF_X1 \buffer_reg[5][3][2][15]  (.D(\input_filter[3][2] [15]), .CK(n_55_7), 
      .Q(\buffer[5][3][2] [15]), .QN());
   DFF_X1 \buffer_reg[5][3][2][14]  (.D(\input_filter[3][2] [14]), .CK(n_55_7), 
      .Q(\buffer[5][3][2] [14]), .QN());
   DFF_X1 \buffer_reg[5][3][2][13]  (.D(\input_filter[3][2] [13]), .CK(n_55_7), 
      .Q(\buffer[5][3][2] [13]), .QN());
   DFF_X1 \buffer_reg[5][3][2][12]  (.D(\input_filter[3][2] [12]), .CK(n_55_7), 
      .Q(\buffer[5][3][2] [12]), .QN());
   DFF_X1 \buffer_reg[5][3][2][11]  (.D(\input_filter[3][2] [11]), .CK(n_55_7), 
      .Q(\buffer[5][3][2] [11]), .QN());
   DFF_X1 \buffer_reg[5][3][2][10]  (.D(\input_filter[3][2] [10]), .CK(n_55_7), 
      .Q(\buffer[5][3][2] [10]), .QN());
   DFF_X1 \buffer_reg[5][3][2][9]  (.D(\input_filter[3][2] [9]), .CK(n_55_7), 
      .Q(\buffer[5][3][2] [9]), .QN());
   DFF_X1 \buffer_reg[5][3][2][8]  (.D(\input_filter[3][2] [8]), .CK(n_55_7), 
      .Q(\buffer[5][3][2] [8]), .QN());
   DFF_X1 \buffer_reg[5][3][2][7]  (.D(\input_filter[3][2] [7]), .CK(n_55_7), 
      .Q(\buffer[5][3][2] [7]), .QN());
   DFF_X1 \buffer_reg[5][3][2][6]  (.D(\input_filter[3][2] [6]), .CK(n_55_7), 
      .Q(\buffer[5][3][2] [6]), .QN());
   DFF_X1 \buffer_reg[5][3][2][5]  (.D(\input_filter[3][2] [5]), .CK(n_55_7), 
      .Q(\buffer[5][3][2] [5]), .QN());
   DFF_X1 \buffer_reg[5][3][2][4]  (.D(\input_filter[3][2] [4]), .CK(n_55_7), 
      .Q(\buffer[5][3][2] [4]), .QN());
   DFF_X1 \buffer_reg[5][3][2][3]  (.D(\input_filter[3][2] [3]), .CK(n_55_7), 
      .Q(\buffer[5][3][2] [3]), .QN());
   DFF_X1 \buffer_reg[5][3][2][2]  (.D(\input_filter[3][2] [2]), .CK(n_55_7), 
      .Q(\buffer[5][3][2] [2]), .QN());
   DFF_X1 \buffer_reg[5][3][2][1]  (.D(\input_filter[3][2] [1]), .CK(n_55_7), 
      .Q(\buffer[5][3][2] [1]), .QN());
   DFF_X1 \buffer_reg[5][3][2][0]  (.D(\input_filter[3][2] [0]), .CK(n_55_7), 
      .Q(\buffer[5][3][2] [0]), .QN());
   DFF_X1 \buffer_reg[4][3][2][15]  (.D(\input_filter[3][2] [15]), .CK(n_55_8), 
      .Q(\buffer[4][3][2] [15]), .QN());
   DFF_X1 \buffer_reg[4][3][2][14]  (.D(\input_filter[3][2] [14]), .CK(n_55_8), 
      .Q(\buffer[4][3][2] [14]), .QN());
   DFF_X1 \buffer_reg[4][3][2][13]  (.D(\input_filter[3][2] [13]), .CK(n_55_8), 
      .Q(\buffer[4][3][2] [13]), .QN());
   DFF_X1 \buffer_reg[4][3][2][12]  (.D(\input_filter[3][2] [12]), .CK(n_55_8), 
      .Q(\buffer[4][3][2] [12]), .QN());
   DFF_X1 \buffer_reg[4][3][2][11]  (.D(\input_filter[3][2] [11]), .CK(n_55_8), 
      .Q(\buffer[4][3][2] [11]), .QN());
   DFF_X1 \buffer_reg[4][3][2][10]  (.D(\input_filter[3][2] [10]), .CK(n_55_8), 
      .Q(\buffer[4][3][2] [10]), .QN());
   DFF_X1 \buffer_reg[4][3][2][9]  (.D(\input_filter[3][2] [9]), .CK(n_55_8), 
      .Q(\buffer[4][3][2] [9]), .QN());
   DFF_X1 \buffer_reg[4][3][2][8]  (.D(\input_filter[3][2] [8]), .CK(n_55_8), 
      .Q(\buffer[4][3][2] [8]), .QN());
   DFF_X1 \buffer_reg[4][3][2][7]  (.D(\input_filter[3][2] [7]), .CK(n_55_8), 
      .Q(\buffer[4][3][2] [7]), .QN());
   DFF_X1 \buffer_reg[4][3][2][6]  (.D(\input_filter[3][2] [6]), .CK(n_55_8), 
      .Q(\buffer[4][3][2] [6]), .QN());
   DFF_X1 \buffer_reg[4][3][2][5]  (.D(\input_filter[3][2] [5]), .CK(n_55_8), 
      .Q(\buffer[4][3][2] [5]), .QN());
   DFF_X1 \buffer_reg[4][3][2][4]  (.D(\input_filter[3][2] [4]), .CK(n_55_8), 
      .Q(\buffer[4][3][2] [4]), .QN());
   DFF_X1 \buffer_reg[4][3][2][3]  (.D(\input_filter[3][2] [3]), .CK(n_55_8), 
      .Q(\buffer[4][3][2] [3]), .QN());
   DFF_X1 \buffer_reg[4][3][2][2]  (.D(\input_filter[3][2] [2]), .CK(n_55_8), 
      .Q(\buffer[4][3][2] [2]), .QN());
   DFF_X1 \buffer_reg[4][3][2][1]  (.D(\input_filter[3][2] [1]), .CK(n_55_8), 
      .Q(\buffer[4][3][2] [1]), .QN());
   DFF_X1 \buffer_reg[4][3][2][0]  (.D(\input_filter[3][2] [0]), .CK(n_55_8), 
      .Q(\buffer[4][3][2] [0]), .QN());
   DFF_X1 \buffer_reg[3][3][2][15]  (.D(\input_filter[3][2] [15]), .CK(n_55_9), 
      .Q(\buffer[3][3][2] [15]), .QN());
   DFF_X1 \buffer_reg[3][3][2][14]  (.D(\input_filter[3][2] [14]), .CK(n_55_9), 
      .Q(\buffer[3][3][2] [14]), .QN());
   DFF_X1 \buffer_reg[3][3][2][13]  (.D(\input_filter[3][2] [13]), .CK(n_55_9), 
      .Q(\buffer[3][3][2] [13]), .QN());
   DFF_X1 \buffer_reg[3][3][2][12]  (.D(\input_filter[3][2] [12]), .CK(n_55_9), 
      .Q(\buffer[3][3][2] [12]), .QN());
   DFF_X1 \buffer_reg[3][3][2][11]  (.D(\input_filter[3][2] [11]), .CK(n_55_9), 
      .Q(\buffer[3][3][2] [11]), .QN());
   DFF_X1 \buffer_reg[3][3][2][10]  (.D(\input_filter[3][2] [10]), .CK(n_55_9), 
      .Q(\buffer[3][3][2] [10]), .QN());
   DFF_X1 \buffer_reg[3][3][2][9]  (.D(\input_filter[3][2] [9]), .CK(n_55_9), 
      .Q(\buffer[3][3][2] [9]), .QN());
   DFF_X1 \buffer_reg[3][3][2][8]  (.D(\input_filter[3][2] [8]), .CK(n_55_9), 
      .Q(\buffer[3][3][2] [8]), .QN());
   DFF_X1 \buffer_reg[3][3][2][7]  (.D(\input_filter[3][2] [7]), .CK(n_55_9), 
      .Q(\buffer[3][3][2] [7]), .QN());
   DFF_X1 \buffer_reg[3][3][2][6]  (.D(\input_filter[3][2] [6]), .CK(n_55_9), 
      .Q(\buffer[3][3][2] [6]), .QN());
   DFF_X1 \buffer_reg[3][3][2][5]  (.D(\input_filter[3][2] [5]), .CK(n_55_9), 
      .Q(\buffer[3][3][2] [5]), .QN());
   DFF_X1 \buffer_reg[3][3][2][4]  (.D(\input_filter[3][2] [4]), .CK(n_55_9), 
      .Q(\buffer[3][3][2] [4]), .QN());
   DFF_X1 \buffer_reg[3][3][2][3]  (.D(\input_filter[3][2] [3]), .CK(n_55_9), 
      .Q(\buffer[3][3][2] [3]), .QN());
   DFF_X1 \buffer_reg[3][3][2][2]  (.D(\input_filter[3][2] [2]), .CK(n_55_9), 
      .Q(\buffer[3][3][2] [2]), .QN());
   DFF_X1 \buffer_reg[3][3][2][1]  (.D(\input_filter[3][2] [1]), .CK(n_55_9), 
      .Q(\buffer[3][3][2] [1]), .QN());
   DFF_X1 \buffer_reg[3][3][2][0]  (.D(\input_filter[3][2] [0]), .CK(n_55_9), 
      .Q(\buffer[3][3][2] [0]), .QN());
   DFF_X1 \buffer_reg[2][3][2][15]  (.D(\input_filter[3][2] [15]), .CK(n_55_10), 
      .Q(\buffer[2][3][2] [15]), .QN());
   DFF_X1 \buffer_reg[2][3][2][14]  (.D(\input_filter[3][2] [14]), .CK(n_55_10), 
      .Q(\buffer[2][3][2] [14]), .QN());
   DFF_X1 \buffer_reg[2][3][2][13]  (.D(\input_filter[3][2] [13]), .CK(n_55_10), 
      .Q(\buffer[2][3][2] [13]), .QN());
   DFF_X1 \buffer_reg[2][3][2][12]  (.D(\input_filter[3][2] [12]), .CK(n_55_10), 
      .Q(\buffer[2][3][2] [12]), .QN());
   DFF_X1 \buffer_reg[2][3][2][11]  (.D(\input_filter[3][2] [11]), .CK(n_55_10), 
      .Q(\buffer[2][3][2] [11]), .QN());
   DFF_X1 \buffer_reg[2][3][2][10]  (.D(\input_filter[3][2] [10]), .CK(n_55_10), 
      .Q(\buffer[2][3][2] [10]), .QN());
   DFF_X1 \buffer_reg[2][3][2][9]  (.D(\input_filter[3][2] [9]), .CK(n_55_10), 
      .Q(\buffer[2][3][2] [9]), .QN());
   DFF_X1 \buffer_reg[2][3][2][8]  (.D(\input_filter[3][2] [8]), .CK(n_55_10), 
      .Q(\buffer[2][3][2] [8]), .QN());
   DFF_X1 \buffer_reg[2][3][2][7]  (.D(\input_filter[3][2] [7]), .CK(n_55_10), 
      .Q(\buffer[2][3][2] [7]), .QN());
   DFF_X1 \buffer_reg[2][3][2][6]  (.D(\input_filter[3][2] [6]), .CK(n_55_10), 
      .Q(\buffer[2][3][2] [6]), .QN());
   DFF_X1 \buffer_reg[2][3][2][5]  (.D(\input_filter[3][2] [5]), .CK(n_55_10), 
      .Q(\buffer[2][3][2] [5]), .QN());
   DFF_X1 \buffer_reg[2][3][2][4]  (.D(\input_filter[3][2] [4]), .CK(n_55_10), 
      .Q(\buffer[2][3][2] [4]), .QN());
   DFF_X1 \buffer_reg[2][3][2][3]  (.D(\input_filter[3][2] [3]), .CK(n_55_10), 
      .Q(\buffer[2][3][2] [3]), .QN());
   DFF_X1 \buffer_reg[2][3][2][2]  (.D(\input_filter[3][2] [2]), .CK(n_55_10), 
      .Q(\buffer[2][3][2] [2]), .QN());
   DFF_X1 \buffer_reg[2][3][2][1]  (.D(\input_filter[3][2] [1]), .CK(n_55_10), 
      .Q(\buffer[2][3][2] [1]), .QN());
   DFF_X1 \buffer_reg[2][3][2][0]  (.D(\input_filter[3][2] [0]), .CK(n_55_10), 
      .Q(\buffer[2][3][2] [0]), .QN());
   DFF_X1 \buffer_reg[1][3][2][15]  (.D(\input_filter[3][2] [15]), .CK(n_55_11), 
      .Q(\buffer[1][3][2] [15]), .QN());
   DFF_X1 \buffer_reg[1][3][2][14]  (.D(\input_filter[3][2] [14]), .CK(n_55_11), 
      .Q(\buffer[1][3][2] [14]), .QN());
   DFF_X1 \buffer_reg[1][3][2][13]  (.D(\input_filter[3][2] [13]), .CK(n_55_11), 
      .Q(\buffer[1][3][2] [13]), .QN());
   DFF_X1 \buffer_reg[1][3][2][12]  (.D(\input_filter[3][2] [12]), .CK(n_55_11), 
      .Q(\buffer[1][3][2] [12]), .QN());
   DFF_X1 \buffer_reg[1][3][2][11]  (.D(\input_filter[3][2] [11]), .CK(n_55_11), 
      .Q(\buffer[1][3][2] [11]), .QN());
   DFF_X1 \buffer_reg[1][3][2][10]  (.D(\input_filter[3][2] [10]), .CK(n_55_11), 
      .Q(\buffer[1][3][2] [10]), .QN());
   DFF_X1 \buffer_reg[1][3][2][9]  (.D(\input_filter[3][2] [9]), .CK(n_55_11), 
      .Q(\buffer[1][3][2] [9]), .QN());
   DFF_X1 \buffer_reg[1][3][2][8]  (.D(\input_filter[3][2] [8]), .CK(n_55_11), 
      .Q(\buffer[1][3][2] [8]), .QN());
   DFF_X1 \buffer_reg[1][3][2][7]  (.D(\input_filter[3][2] [7]), .CK(n_55_11), 
      .Q(\buffer[1][3][2] [7]), .QN());
   DFF_X1 \buffer_reg[1][3][2][6]  (.D(\input_filter[3][2] [6]), .CK(n_55_11), 
      .Q(\buffer[1][3][2] [6]), .QN());
   DFF_X1 \buffer_reg[1][3][2][5]  (.D(\input_filter[3][2] [5]), .CK(n_55_11), 
      .Q(\buffer[1][3][2] [5]), .QN());
   DFF_X1 \buffer_reg[1][3][2][4]  (.D(\input_filter[3][2] [4]), .CK(n_55_11), 
      .Q(\buffer[1][3][2] [4]), .QN());
   DFF_X1 \buffer_reg[1][3][2][3]  (.D(\input_filter[3][2] [3]), .CK(n_55_11), 
      .Q(\buffer[1][3][2] [3]), .QN());
   DFF_X1 \buffer_reg[1][3][2][2]  (.D(\input_filter[3][2] [2]), .CK(n_55_11), 
      .Q(\buffer[1][3][2] [2]), .QN());
   DFF_X1 \buffer_reg[1][3][2][1]  (.D(\input_filter[3][2] [1]), .CK(n_55_11), 
      .Q(\buffer[1][3][2] [1]), .QN());
   DFF_X1 \buffer_reg[1][3][2][0]  (.D(\input_filter[3][2] [0]), .CK(n_55_11), 
      .Q(\buffer[1][3][2] [0]), .QN());
   DFF_X1 \buffer_reg[0][3][2][15]  (.D(\input_filter[3][2] [15]), .CK(n_55_12), 
      .Q(\buffer[0][3][2] [15]), .QN());
   DFF_X1 \buffer_reg[0][3][2][14]  (.D(\input_filter[3][2] [14]), .CK(n_55_12), 
      .Q(\buffer[0][3][2] [14]), .QN());
   DFF_X1 \buffer_reg[0][3][2][13]  (.D(\input_filter[3][2] [13]), .CK(n_55_12), 
      .Q(\buffer[0][3][2] [13]), .QN());
   DFF_X1 \buffer_reg[0][3][2][12]  (.D(\input_filter[3][2] [12]), .CK(n_55_12), 
      .Q(\buffer[0][3][2] [12]), .QN());
   DFF_X1 \buffer_reg[0][3][2][11]  (.D(\input_filter[3][2] [11]), .CK(n_55_12), 
      .Q(\buffer[0][3][2] [11]), .QN());
   DFF_X1 \buffer_reg[0][3][2][10]  (.D(\input_filter[3][2] [10]), .CK(n_55_12), 
      .Q(\buffer[0][3][2] [10]), .QN());
   DFF_X1 \buffer_reg[0][3][2][9]  (.D(\input_filter[3][2] [9]), .CK(n_55_12), 
      .Q(\buffer[0][3][2] [9]), .QN());
   DFF_X1 \buffer_reg[0][3][2][8]  (.D(\input_filter[3][2] [8]), .CK(n_55_12), 
      .Q(\buffer[0][3][2] [8]), .QN());
   DFF_X1 \buffer_reg[0][3][2][7]  (.D(\input_filter[3][2] [7]), .CK(n_55_12), 
      .Q(\buffer[0][3][2] [7]), .QN());
   DFF_X1 \buffer_reg[0][3][2][6]  (.D(\input_filter[3][2] [6]), .CK(n_55_12), 
      .Q(\buffer[0][3][2] [6]), .QN());
   DFF_X1 \buffer_reg[0][3][2][5]  (.D(\input_filter[3][2] [5]), .CK(n_55_12), 
      .Q(\buffer[0][3][2] [5]), .QN());
   DFF_X1 \buffer_reg[0][3][2][4]  (.D(\input_filter[3][2] [4]), .CK(n_55_12), 
      .Q(\buffer[0][3][2] [4]), .QN());
   DFF_X1 \buffer_reg[0][3][2][3]  (.D(\input_filter[3][2] [3]), .CK(n_55_12), 
      .Q(\buffer[0][3][2] [3]), .QN());
   DFF_X1 \buffer_reg[0][3][2][2]  (.D(\input_filter[3][2] [2]), .CK(n_55_12), 
      .Q(\buffer[0][3][2] [2]), .QN());
   DFF_X1 \buffer_reg[0][3][2][1]  (.D(\input_filter[3][2] [1]), .CK(n_55_12), 
      .Q(\buffer[0][3][2] [1]), .QN());
   DFF_X1 \buffer_reg[0][3][2][0]  (.D(\input_filter[3][2] [0]), .CK(n_55_12), 
      .Q(\buffer[0][3][2] [0]), .QN());
   DFF_X1 \buffer_reg[15][3][1][15]  (.D(\input_filter[3][1] [15]), .CK(n_55_13), 
      .Q(\buffer[15][3][1] [15]), .QN());
   DFF_X1 \buffer_reg[15][3][1][14]  (.D(\input_filter[3][1] [14]), .CK(n_55_13), 
      .Q(\buffer[15][3][1] [14]), .QN());
   DFF_X1 \buffer_reg[15][3][1][13]  (.D(\input_filter[3][1] [13]), .CK(n_55_13), 
      .Q(\buffer[15][3][1] [13]), .QN());
   DFF_X1 \buffer_reg[15][3][1][12]  (.D(\input_filter[3][1] [12]), .CK(n_55_13), 
      .Q(\buffer[15][3][1] [12]), .QN());
   DFF_X1 \buffer_reg[15][3][1][11]  (.D(\input_filter[3][1] [11]), .CK(n_55_13), 
      .Q(\buffer[15][3][1] [11]), .QN());
   DFF_X1 \buffer_reg[15][3][1][10]  (.D(\input_filter[3][1] [10]), .CK(n_55_13), 
      .Q(\buffer[15][3][1] [10]), .QN());
   DFF_X1 \buffer_reg[15][3][1][9]  (.D(\input_filter[3][1] [9]), .CK(n_55_13), 
      .Q(\buffer[15][3][1] [9]), .QN());
   DFF_X1 \buffer_reg[15][3][1][8]  (.D(\input_filter[3][1] [8]), .CK(n_55_13), 
      .Q(\buffer[15][3][1] [8]), .QN());
   DFF_X1 \buffer_reg[15][3][1][7]  (.D(\input_filter[3][1] [7]), .CK(n_55_13), 
      .Q(\buffer[15][3][1] [7]), .QN());
   DFF_X1 \buffer_reg[15][3][1][6]  (.D(\input_filter[3][1] [6]), .CK(n_55_13), 
      .Q(\buffer[15][3][1] [6]), .QN());
   DFF_X1 \buffer_reg[15][3][1][5]  (.D(\input_filter[3][1] [5]), .CK(n_55_13), 
      .Q(\buffer[15][3][1] [5]), .QN());
   DFF_X1 \buffer_reg[15][3][1][4]  (.D(\input_filter[3][1] [4]), .CK(n_55_13), 
      .Q(\buffer[15][3][1] [4]), .QN());
   DFF_X1 \buffer_reg[15][3][1][3]  (.D(\input_filter[3][1] [3]), .CK(n_55_13), 
      .Q(\buffer[15][3][1] [3]), .QN());
   DFF_X1 \buffer_reg[15][3][1][2]  (.D(\input_filter[3][1] [2]), .CK(n_55_13), 
      .Q(\buffer[15][3][1] [2]), .QN());
   DFF_X1 \buffer_reg[15][3][1][1]  (.D(\input_filter[3][1] [1]), .CK(n_55_13), 
      .Q(\buffer[15][3][1] [1]), .QN());
   DFF_X1 \buffer_reg[15][3][1][0]  (.D(\input_filter[3][1] [0]), .CK(n_55_13), 
      .Q(\buffer[15][3][1] [0]), .QN());
   DFF_X1 \buffer_reg[14][3][1][15]  (.D(\input_filter[3][1] [15]), .CK(n_55_14), 
      .Q(\buffer[14][3][1] [15]), .QN());
   DFF_X1 \buffer_reg[14][3][1][14]  (.D(\input_filter[3][1] [14]), .CK(n_55_14), 
      .Q(\buffer[14][3][1] [14]), .QN());
   DFF_X1 \buffer_reg[14][3][1][13]  (.D(\input_filter[3][1] [13]), .CK(n_55_14), 
      .Q(\buffer[14][3][1] [13]), .QN());
   DFF_X1 \buffer_reg[14][3][1][12]  (.D(\input_filter[3][1] [12]), .CK(n_55_14), 
      .Q(\buffer[14][3][1] [12]), .QN());
   DFF_X1 \buffer_reg[14][3][1][11]  (.D(\input_filter[3][1] [11]), .CK(n_55_14), 
      .Q(\buffer[14][3][1] [11]), .QN());
   DFF_X1 \buffer_reg[14][3][1][10]  (.D(\input_filter[3][1] [10]), .CK(n_55_14), 
      .Q(\buffer[14][3][1] [10]), .QN());
   DFF_X1 \buffer_reg[14][3][1][9]  (.D(\input_filter[3][1] [9]), .CK(n_55_14), 
      .Q(\buffer[14][3][1] [9]), .QN());
   DFF_X1 \buffer_reg[14][3][1][8]  (.D(\input_filter[3][1] [8]), .CK(n_55_14), 
      .Q(\buffer[14][3][1] [8]), .QN());
   DFF_X1 \buffer_reg[14][3][1][7]  (.D(\input_filter[3][1] [7]), .CK(n_55_14), 
      .Q(\buffer[14][3][1] [7]), .QN());
   DFF_X1 \buffer_reg[14][3][1][6]  (.D(\input_filter[3][1] [6]), .CK(n_55_14), 
      .Q(\buffer[14][3][1] [6]), .QN());
   DFF_X1 \buffer_reg[14][3][1][5]  (.D(\input_filter[3][1] [5]), .CK(n_55_14), 
      .Q(\buffer[14][3][1] [5]), .QN());
   DFF_X1 \buffer_reg[14][3][1][4]  (.D(\input_filter[3][1] [4]), .CK(n_55_14), 
      .Q(\buffer[14][3][1] [4]), .QN());
   DFF_X1 \buffer_reg[14][3][1][3]  (.D(\input_filter[3][1] [3]), .CK(n_55_14), 
      .Q(\buffer[14][3][1] [3]), .QN());
   DFF_X1 \buffer_reg[14][3][1][2]  (.D(\input_filter[3][1] [2]), .CK(n_55_14), 
      .Q(\buffer[14][3][1] [2]), .QN());
   DFF_X1 \buffer_reg[14][3][1][1]  (.D(\input_filter[3][1] [1]), .CK(n_55_14), 
      .Q(\buffer[14][3][1] [1]), .QN());
   DFF_X1 \buffer_reg[14][3][1][0]  (.D(\input_filter[3][1] [0]), .CK(n_55_14), 
      .Q(\buffer[14][3][1] [0]), .QN());
   DFF_X1 \buffer_reg[13][3][1][15]  (.D(\input_filter[3][1] [15]), .CK(n_55_15), 
      .Q(\buffer[13][3][1] [15]), .QN());
   DFF_X1 \buffer_reg[13][3][1][14]  (.D(\input_filter[3][1] [14]), .CK(n_55_15), 
      .Q(\buffer[13][3][1] [14]), .QN());
   DFF_X1 \buffer_reg[13][3][1][13]  (.D(\input_filter[3][1] [13]), .CK(n_55_15), 
      .Q(\buffer[13][3][1] [13]), .QN());
   DFF_X1 \buffer_reg[13][3][1][12]  (.D(\input_filter[3][1] [12]), .CK(n_55_15), 
      .Q(\buffer[13][3][1] [12]), .QN());
   DFF_X1 \buffer_reg[13][3][1][11]  (.D(\input_filter[3][1] [11]), .CK(n_55_15), 
      .Q(\buffer[13][3][1] [11]), .QN());
   DFF_X1 \buffer_reg[13][3][1][10]  (.D(\input_filter[3][1] [10]), .CK(n_55_15), 
      .Q(\buffer[13][3][1] [10]), .QN());
   DFF_X1 \buffer_reg[13][3][1][9]  (.D(\input_filter[3][1] [9]), .CK(n_55_15), 
      .Q(\buffer[13][3][1] [9]), .QN());
   DFF_X1 \buffer_reg[13][3][1][8]  (.D(\input_filter[3][1] [8]), .CK(n_55_15), 
      .Q(\buffer[13][3][1] [8]), .QN());
   DFF_X1 \buffer_reg[13][3][1][7]  (.D(\input_filter[3][1] [7]), .CK(n_55_15), 
      .Q(\buffer[13][3][1] [7]), .QN());
   DFF_X1 \buffer_reg[13][3][1][6]  (.D(\input_filter[3][1] [6]), .CK(n_55_15), 
      .Q(\buffer[13][3][1] [6]), .QN());
   DFF_X1 \buffer_reg[13][3][1][5]  (.D(\input_filter[3][1] [5]), .CK(n_55_15), 
      .Q(\buffer[13][3][1] [5]), .QN());
   DFF_X1 \buffer_reg[13][3][1][4]  (.D(\input_filter[3][1] [4]), .CK(n_55_15), 
      .Q(\buffer[13][3][1] [4]), .QN());
   DFF_X1 \buffer_reg[13][3][1][3]  (.D(\input_filter[3][1] [3]), .CK(n_55_15), 
      .Q(\buffer[13][3][1] [3]), .QN());
   DFF_X1 \buffer_reg[13][3][1][2]  (.D(\input_filter[3][1] [2]), .CK(n_55_15), 
      .Q(\buffer[13][3][1] [2]), .QN());
   DFF_X1 \buffer_reg[13][3][1][1]  (.D(\input_filter[3][1] [1]), .CK(n_55_15), 
      .Q(\buffer[13][3][1] [1]), .QN());
   DFF_X1 \buffer_reg[13][3][1][0]  (.D(\input_filter[3][1] [0]), .CK(n_55_15), 
      .Q(\buffer[13][3][1] [0]), .QN());
   DFF_X1 \buffer_reg[12][3][1][15]  (.D(\input_filter[3][1] [15]), .CK(n_55_0), 
      .Q(\buffer[12][3][1] [15]), .QN());
   DFF_X1 \buffer_reg[12][3][1][14]  (.D(\input_filter[3][1] [14]), .CK(n_55_0), 
      .Q(\buffer[12][3][1] [14]), .QN());
   DFF_X1 \buffer_reg[12][3][1][13]  (.D(\input_filter[3][1] [13]), .CK(n_55_0), 
      .Q(\buffer[12][3][1] [13]), .QN());
   DFF_X1 \buffer_reg[12][3][1][12]  (.D(\input_filter[3][1] [12]), .CK(n_55_0), 
      .Q(\buffer[12][3][1] [12]), .QN());
   DFF_X1 \buffer_reg[12][3][1][11]  (.D(\input_filter[3][1] [11]), .CK(n_55_0), 
      .Q(\buffer[12][3][1] [11]), .QN());
   DFF_X1 \buffer_reg[12][3][1][10]  (.D(\input_filter[3][1] [10]), .CK(n_55_0), 
      .Q(\buffer[12][3][1] [10]), .QN());
   DFF_X1 \buffer_reg[12][3][1][9]  (.D(\input_filter[3][1] [9]), .CK(n_55_0), 
      .Q(\buffer[12][3][1] [9]), .QN());
   DFF_X1 \buffer_reg[12][3][1][8]  (.D(\input_filter[3][1] [8]), .CK(n_55_0), 
      .Q(\buffer[12][3][1] [8]), .QN());
   DFF_X1 \buffer_reg[12][3][1][7]  (.D(\input_filter[3][1] [7]), .CK(n_55_0), 
      .Q(\buffer[12][3][1] [7]), .QN());
   DFF_X1 \buffer_reg[12][3][1][6]  (.D(\input_filter[3][1] [6]), .CK(n_55_0), 
      .Q(\buffer[12][3][1] [6]), .QN());
   DFF_X1 \buffer_reg[12][3][1][5]  (.D(\input_filter[3][1] [5]), .CK(n_55_0), 
      .Q(\buffer[12][3][1] [5]), .QN());
   DFF_X1 \buffer_reg[12][3][1][4]  (.D(\input_filter[3][1] [4]), .CK(n_55_0), 
      .Q(\buffer[12][3][1] [4]), .QN());
   DFF_X1 \buffer_reg[12][3][1][3]  (.D(\input_filter[3][1] [3]), .CK(n_55_0), 
      .Q(\buffer[12][3][1] [3]), .QN());
   DFF_X1 \buffer_reg[12][3][1][2]  (.D(\input_filter[3][1] [2]), .CK(n_55_0), 
      .Q(\buffer[12][3][1] [2]), .QN());
   DFF_X1 \buffer_reg[12][3][1][1]  (.D(\input_filter[3][1] [1]), .CK(n_55_0), 
      .Q(\buffer[12][3][1] [1]), .QN());
   DFF_X1 \buffer_reg[12][3][1][0]  (.D(\input_filter[3][1] [0]), .CK(n_55_0), 
      .Q(\buffer[12][3][1] [0]), .QN());
   DFF_X1 \buffer_reg[11][3][1][15]  (.D(\input_filter[3][1] [15]), .CK(n_55_1), 
      .Q(\buffer[11][3][1] [15]), .QN());
   DFF_X1 \buffer_reg[11][3][1][14]  (.D(\input_filter[3][1] [14]), .CK(n_55_1), 
      .Q(\buffer[11][3][1] [14]), .QN());
   DFF_X1 \buffer_reg[11][3][1][13]  (.D(\input_filter[3][1] [13]), .CK(n_55_1), 
      .Q(\buffer[11][3][1] [13]), .QN());
   DFF_X1 \buffer_reg[11][3][1][12]  (.D(\input_filter[3][1] [12]), .CK(n_55_1), 
      .Q(\buffer[11][3][1] [12]), .QN());
   DFF_X1 \buffer_reg[11][3][1][11]  (.D(\input_filter[3][1] [11]), .CK(n_55_1), 
      .Q(\buffer[11][3][1] [11]), .QN());
   DFF_X1 \buffer_reg[11][3][1][10]  (.D(\input_filter[3][1] [10]), .CK(n_55_1), 
      .Q(\buffer[11][3][1] [10]), .QN());
   DFF_X1 \buffer_reg[11][3][1][9]  (.D(\input_filter[3][1] [9]), .CK(n_55_1), 
      .Q(\buffer[11][3][1] [9]), .QN());
   DFF_X1 \buffer_reg[11][3][1][8]  (.D(\input_filter[3][1] [8]), .CK(n_55_1), 
      .Q(\buffer[11][3][1] [8]), .QN());
   DFF_X1 \buffer_reg[11][3][1][7]  (.D(\input_filter[3][1] [7]), .CK(n_55_1), 
      .Q(\buffer[11][3][1] [7]), .QN());
   DFF_X1 \buffer_reg[11][3][1][6]  (.D(\input_filter[3][1] [6]), .CK(n_55_1), 
      .Q(\buffer[11][3][1] [6]), .QN());
   DFF_X1 \buffer_reg[11][3][1][5]  (.D(\input_filter[3][1] [5]), .CK(n_55_1), 
      .Q(\buffer[11][3][1] [5]), .QN());
   DFF_X1 \buffer_reg[11][3][1][4]  (.D(\input_filter[3][1] [4]), .CK(n_55_1), 
      .Q(\buffer[11][3][1] [4]), .QN());
   DFF_X1 \buffer_reg[11][3][1][3]  (.D(\input_filter[3][1] [3]), .CK(n_55_1), 
      .Q(\buffer[11][3][1] [3]), .QN());
   DFF_X1 \buffer_reg[11][3][1][2]  (.D(\input_filter[3][1] [2]), .CK(n_55_1), 
      .Q(\buffer[11][3][1] [2]), .QN());
   DFF_X1 \buffer_reg[11][3][1][1]  (.D(\input_filter[3][1] [1]), .CK(n_55_1), 
      .Q(\buffer[11][3][1] [1]), .QN());
   DFF_X1 \buffer_reg[11][3][1][0]  (.D(\input_filter[3][1] [0]), .CK(n_55_1), 
      .Q(\buffer[11][3][1] [0]), .QN());
   DFF_X1 \buffer_reg[10][3][1][15]  (.D(\input_filter[3][1] [15]), .CK(n_55_2), 
      .Q(\buffer[10][3][1] [15]), .QN());
   DFF_X1 \buffer_reg[10][3][1][14]  (.D(\input_filter[3][1] [14]), .CK(n_55_2), 
      .Q(\buffer[10][3][1] [14]), .QN());
   DFF_X1 \buffer_reg[10][3][1][13]  (.D(\input_filter[3][1] [13]), .CK(n_55_2), 
      .Q(\buffer[10][3][1] [13]), .QN());
   DFF_X1 \buffer_reg[10][3][1][12]  (.D(\input_filter[3][1] [12]), .CK(n_55_2), 
      .Q(\buffer[10][3][1] [12]), .QN());
   DFF_X1 \buffer_reg[10][3][1][11]  (.D(\input_filter[3][1] [11]), .CK(n_55_2), 
      .Q(\buffer[10][3][1] [11]), .QN());
   DFF_X1 \buffer_reg[10][3][1][10]  (.D(\input_filter[3][1] [10]), .CK(n_55_2), 
      .Q(\buffer[10][3][1] [10]), .QN());
   DFF_X1 \buffer_reg[10][3][1][9]  (.D(\input_filter[3][1] [9]), .CK(n_55_2), 
      .Q(\buffer[10][3][1] [9]), .QN());
   DFF_X1 \buffer_reg[10][3][1][8]  (.D(\input_filter[3][1] [8]), .CK(n_55_2), 
      .Q(\buffer[10][3][1] [8]), .QN());
   DFF_X1 \buffer_reg[10][3][1][7]  (.D(\input_filter[3][1] [7]), .CK(n_55_2), 
      .Q(\buffer[10][3][1] [7]), .QN());
   DFF_X1 \buffer_reg[10][3][1][6]  (.D(\input_filter[3][1] [6]), .CK(n_55_2), 
      .Q(\buffer[10][3][1] [6]), .QN());
   DFF_X1 \buffer_reg[10][3][1][5]  (.D(\input_filter[3][1] [5]), .CK(n_55_2), 
      .Q(\buffer[10][3][1] [5]), .QN());
   DFF_X1 \buffer_reg[10][3][1][4]  (.D(\input_filter[3][1] [4]), .CK(n_55_2), 
      .Q(\buffer[10][3][1] [4]), .QN());
   DFF_X1 \buffer_reg[10][3][1][3]  (.D(\input_filter[3][1] [3]), .CK(n_55_2), 
      .Q(\buffer[10][3][1] [3]), .QN());
   DFF_X1 \buffer_reg[10][3][1][2]  (.D(\input_filter[3][1] [2]), .CK(n_55_2), 
      .Q(\buffer[10][3][1] [2]), .QN());
   DFF_X1 \buffer_reg[10][3][1][1]  (.D(\input_filter[3][1] [1]), .CK(n_55_2), 
      .Q(\buffer[10][3][1] [1]), .QN());
   DFF_X1 \buffer_reg[10][3][1][0]  (.D(\input_filter[3][1] [0]), .CK(n_55_2), 
      .Q(\buffer[10][3][1] [0]), .QN());
   DFF_X1 \buffer_reg[9][3][1][15]  (.D(\input_filter[3][1] [15]), .CK(n_55_3), 
      .Q(\buffer[9][3][1] [15]), .QN());
   DFF_X1 \buffer_reg[9][3][1][14]  (.D(\input_filter[3][1] [14]), .CK(n_55_3), 
      .Q(\buffer[9][3][1] [14]), .QN());
   DFF_X1 \buffer_reg[9][3][1][13]  (.D(\input_filter[3][1] [13]), .CK(n_55_3), 
      .Q(\buffer[9][3][1] [13]), .QN());
   DFF_X1 \buffer_reg[9][3][1][12]  (.D(\input_filter[3][1] [12]), .CK(n_55_3), 
      .Q(\buffer[9][3][1] [12]), .QN());
   DFF_X1 \buffer_reg[9][3][1][11]  (.D(\input_filter[3][1] [11]), .CK(n_55_3), 
      .Q(\buffer[9][3][1] [11]), .QN());
   DFF_X1 \buffer_reg[9][3][1][10]  (.D(\input_filter[3][1] [10]), .CK(n_55_3), 
      .Q(\buffer[9][3][1] [10]), .QN());
   DFF_X1 \buffer_reg[9][3][1][9]  (.D(\input_filter[3][1] [9]), .CK(n_55_3), 
      .Q(\buffer[9][3][1] [9]), .QN());
   DFF_X1 \buffer_reg[9][3][1][8]  (.D(\input_filter[3][1] [8]), .CK(n_55_3), 
      .Q(\buffer[9][3][1] [8]), .QN());
   DFF_X1 \buffer_reg[9][3][1][7]  (.D(\input_filter[3][1] [7]), .CK(n_55_3), 
      .Q(\buffer[9][3][1] [7]), .QN());
   DFF_X1 \buffer_reg[9][3][1][6]  (.D(\input_filter[3][1] [6]), .CK(n_55_3), 
      .Q(\buffer[9][3][1] [6]), .QN());
   DFF_X1 \buffer_reg[9][3][1][5]  (.D(\input_filter[3][1] [5]), .CK(n_55_3), 
      .Q(\buffer[9][3][1] [5]), .QN());
   DFF_X1 \buffer_reg[9][3][1][4]  (.D(\input_filter[3][1] [4]), .CK(n_55_3), 
      .Q(\buffer[9][3][1] [4]), .QN());
   DFF_X1 \buffer_reg[9][3][1][3]  (.D(\input_filter[3][1] [3]), .CK(n_55_3), 
      .Q(\buffer[9][3][1] [3]), .QN());
   DFF_X1 \buffer_reg[9][3][1][2]  (.D(\input_filter[3][1] [2]), .CK(n_55_3), 
      .Q(\buffer[9][3][1] [2]), .QN());
   DFF_X1 \buffer_reg[9][3][1][1]  (.D(\input_filter[3][1] [1]), .CK(n_55_3), 
      .Q(\buffer[9][3][1] [1]), .QN());
   DFF_X1 \buffer_reg[9][3][1][0]  (.D(\input_filter[3][1] [0]), .CK(n_55_3), 
      .Q(\buffer[9][3][1] [0]), .QN());
   DFF_X1 \buffer_reg[8][3][1][15]  (.D(\input_filter[3][1] [15]), .CK(n_55_4), 
      .Q(\buffer[8][3][1] [15]), .QN());
   DFF_X1 \buffer_reg[8][3][1][14]  (.D(\input_filter[3][1] [14]), .CK(n_55_4), 
      .Q(\buffer[8][3][1] [14]), .QN());
   DFF_X1 \buffer_reg[8][3][1][13]  (.D(\input_filter[3][1] [13]), .CK(n_55_4), 
      .Q(\buffer[8][3][1] [13]), .QN());
   DFF_X1 \buffer_reg[8][3][1][12]  (.D(\input_filter[3][1] [12]), .CK(n_55_4), 
      .Q(\buffer[8][3][1] [12]), .QN());
   DFF_X1 \buffer_reg[8][3][1][11]  (.D(\input_filter[3][1] [11]), .CK(n_55_4), 
      .Q(\buffer[8][3][1] [11]), .QN());
   DFF_X1 \buffer_reg[8][3][1][10]  (.D(\input_filter[3][1] [10]), .CK(n_55_4), 
      .Q(\buffer[8][3][1] [10]), .QN());
   DFF_X1 \buffer_reg[8][3][1][9]  (.D(\input_filter[3][1] [9]), .CK(n_55_4), 
      .Q(\buffer[8][3][1] [9]), .QN());
   DFF_X1 \buffer_reg[8][3][1][8]  (.D(\input_filter[3][1] [8]), .CK(n_55_4), 
      .Q(\buffer[8][3][1] [8]), .QN());
   DFF_X1 \buffer_reg[8][3][1][7]  (.D(\input_filter[3][1] [7]), .CK(n_55_4), 
      .Q(\buffer[8][3][1] [7]), .QN());
   DFF_X1 \buffer_reg[8][3][1][6]  (.D(\input_filter[3][1] [6]), .CK(n_55_4), 
      .Q(\buffer[8][3][1] [6]), .QN());
   DFF_X1 \buffer_reg[8][3][1][5]  (.D(\input_filter[3][1] [5]), .CK(n_55_4), 
      .Q(\buffer[8][3][1] [5]), .QN());
   DFF_X1 \buffer_reg[8][3][1][4]  (.D(\input_filter[3][1] [4]), .CK(n_55_4), 
      .Q(\buffer[8][3][1] [4]), .QN());
   DFF_X1 \buffer_reg[8][3][1][3]  (.D(\input_filter[3][1] [3]), .CK(n_55_4), 
      .Q(\buffer[8][3][1] [3]), .QN());
   DFF_X1 \buffer_reg[8][3][1][2]  (.D(\input_filter[3][1] [2]), .CK(n_55_4), 
      .Q(\buffer[8][3][1] [2]), .QN());
   DFF_X1 \buffer_reg[8][3][1][1]  (.D(\input_filter[3][1] [1]), .CK(n_55_4), 
      .Q(\buffer[8][3][1] [1]), .QN());
   DFF_X1 \buffer_reg[8][3][1][0]  (.D(\input_filter[3][1] [0]), .CK(n_55_4), 
      .Q(\buffer[8][3][1] [0]), .QN());
   DFF_X1 \buffer_reg[7][3][1][15]  (.D(\input_filter[3][1] [15]), .CK(n_55_5), 
      .Q(\buffer[7][3][1] [15]), .QN());
   DFF_X1 \buffer_reg[7][3][1][14]  (.D(\input_filter[3][1] [14]), .CK(n_55_5), 
      .Q(\buffer[7][3][1] [14]), .QN());
   DFF_X1 \buffer_reg[7][3][1][13]  (.D(\input_filter[3][1] [13]), .CK(n_55_5), 
      .Q(\buffer[7][3][1] [13]), .QN());
   DFF_X1 \buffer_reg[7][3][1][12]  (.D(\input_filter[3][1] [12]), .CK(n_55_5), 
      .Q(\buffer[7][3][1] [12]), .QN());
   DFF_X1 \buffer_reg[7][3][1][11]  (.D(\input_filter[3][1] [11]), .CK(n_55_5), 
      .Q(\buffer[7][3][1] [11]), .QN());
   DFF_X1 \buffer_reg[7][3][1][10]  (.D(\input_filter[3][1] [10]), .CK(n_55_5), 
      .Q(\buffer[7][3][1] [10]), .QN());
   DFF_X1 \buffer_reg[7][3][1][9]  (.D(\input_filter[3][1] [9]), .CK(n_55_5), 
      .Q(\buffer[7][3][1] [9]), .QN());
   DFF_X1 \buffer_reg[7][3][1][8]  (.D(\input_filter[3][1] [8]), .CK(n_55_5), 
      .Q(\buffer[7][3][1] [8]), .QN());
   DFF_X1 \buffer_reg[7][3][1][7]  (.D(\input_filter[3][1] [7]), .CK(n_55_5), 
      .Q(\buffer[7][3][1] [7]), .QN());
   DFF_X1 \buffer_reg[7][3][1][6]  (.D(\input_filter[3][1] [6]), .CK(n_55_5), 
      .Q(\buffer[7][3][1] [6]), .QN());
   DFF_X1 \buffer_reg[7][3][1][5]  (.D(\input_filter[3][1] [5]), .CK(n_55_5), 
      .Q(\buffer[7][3][1] [5]), .QN());
   DFF_X1 \buffer_reg[7][3][1][4]  (.D(\input_filter[3][1] [4]), .CK(n_55_5), 
      .Q(\buffer[7][3][1] [4]), .QN());
   DFF_X1 \buffer_reg[7][3][1][3]  (.D(\input_filter[3][1] [3]), .CK(n_55_5), 
      .Q(\buffer[7][3][1] [3]), .QN());
   DFF_X1 \buffer_reg[7][3][1][2]  (.D(\input_filter[3][1] [2]), .CK(n_55_5), 
      .Q(\buffer[7][3][1] [2]), .QN());
   DFF_X1 \buffer_reg[7][3][1][1]  (.D(\input_filter[3][1] [1]), .CK(n_55_5), 
      .Q(\buffer[7][3][1] [1]), .QN());
   DFF_X1 \buffer_reg[7][3][1][0]  (.D(\input_filter[3][1] [0]), .CK(n_55_5), 
      .Q(\buffer[7][3][1] [0]), .QN());
   DFF_X1 \buffer_reg[6][3][1][15]  (.D(\input_filter[3][1] [15]), .CK(n_55_6), 
      .Q(\buffer[6][3][1] [15]), .QN());
   DFF_X1 \buffer_reg[6][3][1][14]  (.D(\input_filter[3][1] [14]), .CK(n_55_6), 
      .Q(\buffer[6][3][1] [14]), .QN());
   DFF_X1 \buffer_reg[6][3][1][13]  (.D(\input_filter[3][1] [13]), .CK(n_55_6), 
      .Q(\buffer[6][3][1] [13]), .QN());
   DFF_X1 \buffer_reg[6][3][1][12]  (.D(\input_filter[3][1] [12]), .CK(n_55_6), 
      .Q(\buffer[6][3][1] [12]), .QN());
   DFF_X1 \buffer_reg[6][3][1][11]  (.D(\input_filter[3][1] [11]), .CK(n_55_6), 
      .Q(\buffer[6][3][1] [11]), .QN());
   DFF_X1 \buffer_reg[6][3][1][10]  (.D(\input_filter[3][1] [10]), .CK(n_55_6), 
      .Q(\buffer[6][3][1] [10]), .QN());
   DFF_X1 \buffer_reg[6][3][1][9]  (.D(\input_filter[3][1] [9]), .CK(n_55_6), 
      .Q(\buffer[6][3][1] [9]), .QN());
   DFF_X1 \buffer_reg[6][3][1][8]  (.D(\input_filter[3][1] [8]), .CK(n_55_6), 
      .Q(\buffer[6][3][1] [8]), .QN());
   DFF_X1 \buffer_reg[6][3][1][7]  (.D(\input_filter[3][1] [7]), .CK(n_55_6), 
      .Q(\buffer[6][3][1] [7]), .QN());
   DFF_X1 \buffer_reg[6][3][1][6]  (.D(\input_filter[3][1] [6]), .CK(n_55_6), 
      .Q(\buffer[6][3][1] [6]), .QN());
   DFF_X1 \buffer_reg[6][3][1][5]  (.D(\input_filter[3][1] [5]), .CK(n_55_6), 
      .Q(\buffer[6][3][1] [5]), .QN());
   DFF_X1 \buffer_reg[6][3][1][4]  (.D(\input_filter[3][1] [4]), .CK(n_55_6), 
      .Q(\buffer[6][3][1] [4]), .QN());
   DFF_X1 \buffer_reg[6][3][1][3]  (.D(\input_filter[3][1] [3]), .CK(n_55_6), 
      .Q(\buffer[6][3][1] [3]), .QN());
   DFF_X1 \buffer_reg[6][3][1][2]  (.D(\input_filter[3][1] [2]), .CK(n_55_6), 
      .Q(\buffer[6][3][1] [2]), .QN());
   DFF_X1 \buffer_reg[6][3][1][1]  (.D(\input_filter[3][1] [1]), .CK(n_55_6), 
      .Q(\buffer[6][3][1] [1]), .QN());
   DFF_X1 \buffer_reg[6][3][1][0]  (.D(\input_filter[3][1] [0]), .CK(n_55_6), 
      .Q(\buffer[6][3][1] [0]), .QN());
   DFF_X1 \buffer_reg[5][3][1][15]  (.D(\input_filter[3][1] [15]), .CK(n_55_7), 
      .Q(\buffer[5][3][1] [15]), .QN());
   DFF_X1 \buffer_reg[5][3][1][14]  (.D(\input_filter[3][1] [14]), .CK(n_55_7), 
      .Q(\buffer[5][3][1] [14]), .QN());
   DFF_X1 \buffer_reg[5][3][1][13]  (.D(\input_filter[3][1] [13]), .CK(n_55_7), 
      .Q(\buffer[5][3][1] [13]), .QN());
   DFF_X1 \buffer_reg[5][3][1][12]  (.D(\input_filter[3][1] [12]), .CK(n_55_7), 
      .Q(\buffer[5][3][1] [12]), .QN());
   DFF_X1 \buffer_reg[5][3][1][11]  (.D(\input_filter[3][1] [11]), .CK(n_55_7), 
      .Q(\buffer[5][3][1] [11]), .QN());
   DFF_X1 \buffer_reg[5][3][1][10]  (.D(\input_filter[3][1] [10]), .CK(n_55_7), 
      .Q(\buffer[5][3][1] [10]), .QN());
   DFF_X1 \buffer_reg[5][3][1][9]  (.D(\input_filter[3][1] [9]), .CK(n_55_7), 
      .Q(\buffer[5][3][1] [9]), .QN());
   DFF_X1 \buffer_reg[5][3][1][8]  (.D(\input_filter[3][1] [8]), .CK(n_55_7), 
      .Q(\buffer[5][3][1] [8]), .QN());
   DFF_X1 \buffer_reg[5][3][1][7]  (.D(\input_filter[3][1] [7]), .CK(n_55_7), 
      .Q(\buffer[5][3][1] [7]), .QN());
   DFF_X1 \buffer_reg[5][3][1][6]  (.D(\input_filter[3][1] [6]), .CK(n_55_7), 
      .Q(\buffer[5][3][1] [6]), .QN());
   DFF_X1 \buffer_reg[5][3][1][5]  (.D(\input_filter[3][1] [5]), .CK(n_55_7), 
      .Q(\buffer[5][3][1] [5]), .QN());
   DFF_X1 \buffer_reg[5][3][1][4]  (.D(\input_filter[3][1] [4]), .CK(n_55_7), 
      .Q(\buffer[5][3][1] [4]), .QN());
   DFF_X1 \buffer_reg[5][3][1][3]  (.D(\input_filter[3][1] [3]), .CK(n_55_7), 
      .Q(\buffer[5][3][1] [3]), .QN());
   DFF_X1 \buffer_reg[5][3][1][2]  (.D(\input_filter[3][1] [2]), .CK(n_55_7), 
      .Q(\buffer[5][3][1] [2]), .QN());
   DFF_X1 \buffer_reg[5][3][1][1]  (.D(\input_filter[3][1] [1]), .CK(n_55_7), 
      .Q(\buffer[5][3][1] [1]), .QN());
   DFF_X1 \buffer_reg[5][3][1][0]  (.D(\input_filter[3][1] [0]), .CK(n_55_7), 
      .Q(\buffer[5][3][1] [0]), .QN());
   DFF_X1 \buffer_reg[4][3][1][15]  (.D(\input_filter[3][1] [15]), .CK(n_55_8), 
      .Q(\buffer[4][3][1] [15]), .QN());
   DFF_X1 \buffer_reg[4][3][1][14]  (.D(\input_filter[3][1] [14]), .CK(n_55_8), 
      .Q(\buffer[4][3][1] [14]), .QN());
   DFF_X1 \buffer_reg[4][3][1][13]  (.D(\input_filter[3][1] [13]), .CK(n_55_8), 
      .Q(\buffer[4][3][1] [13]), .QN());
   DFF_X1 \buffer_reg[4][3][1][12]  (.D(\input_filter[3][1] [12]), .CK(n_55_8), 
      .Q(\buffer[4][3][1] [12]), .QN());
   DFF_X1 \buffer_reg[4][3][1][11]  (.D(\input_filter[3][1] [11]), .CK(n_55_8), 
      .Q(\buffer[4][3][1] [11]), .QN());
   DFF_X1 \buffer_reg[4][3][1][10]  (.D(\input_filter[3][1] [10]), .CK(n_55_8), 
      .Q(\buffer[4][3][1] [10]), .QN());
   DFF_X1 \buffer_reg[4][3][1][9]  (.D(\input_filter[3][1] [9]), .CK(n_55_8), 
      .Q(\buffer[4][3][1] [9]), .QN());
   DFF_X1 \buffer_reg[4][3][1][8]  (.D(\input_filter[3][1] [8]), .CK(n_55_8), 
      .Q(\buffer[4][3][1] [8]), .QN());
   DFF_X1 \buffer_reg[4][3][1][7]  (.D(\input_filter[3][1] [7]), .CK(n_55_8), 
      .Q(\buffer[4][3][1] [7]), .QN());
   DFF_X1 \buffer_reg[4][3][1][6]  (.D(\input_filter[3][1] [6]), .CK(n_55_8), 
      .Q(\buffer[4][3][1] [6]), .QN());
   DFF_X1 \buffer_reg[4][3][1][5]  (.D(\input_filter[3][1] [5]), .CK(n_55_8), 
      .Q(\buffer[4][3][1] [5]), .QN());
   DFF_X1 \buffer_reg[4][3][1][4]  (.D(\input_filter[3][1] [4]), .CK(n_55_8), 
      .Q(\buffer[4][3][1] [4]), .QN());
   DFF_X1 \buffer_reg[4][3][1][3]  (.D(\input_filter[3][1] [3]), .CK(n_55_8), 
      .Q(\buffer[4][3][1] [3]), .QN());
   DFF_X1 \buffer_reg[4][3][1][2]  (.D(\input_filter[3][1] [2]), .CK(n_55_8), 
      .Q(\buffer[4][3][1] [2]), .QN());
   DFF_X1 \buffer_reg[4][3][1][1]  (.D(\input_filter[3][1] [1]), .CK(n_55_8), 
      .Q(\buffer[4][3][1] [1]), .QN());
   DFF_X1 \buffer_reg[4][3][1][0]  (.D(\input_filter[3][1] [0]), .CK(n_55_8), 
      .Q(\buffer[4][3][1] [0]), .QN());
   DFF_X1 \buffer_reg[3][3][1][15]  (.D(\input_filter[3][1] [15]), .CK(n_55_9), 
      .Q(\buffer[3][3][1] [15]), .QN());
   DFF_X1 \buffer_reg[3][3][1][14]  (.D(\input_filter[3][1] [14]), .CK(n_55_9), 
      .Q(\buffer[3][3][1] [14]), .QN());
   DFF_X1 \buffer_reg[3][3][1][13]  (.D(\input_filter[3][1] [13]), .CK(n_55_9), 
      .Q(\buffer[3][3][1] [13]), .QN());
   DFF_X1 \buffer_reg[3][3][1][12]  (.D(\input_filter[3][1] [12]), .CK(n_55_9), 
      .Q(\buffer[3][3][1] [12]), .QN());
   DFF_X1 \buffer_reg[3][3][1][11]  (.D(\input_filter[3][1] [11]), .CK(n_55_9), 
      .Q(\buffer[3][3][1] [11]), .QN());
   DFF_X1 \buffer_reg[3][3][1][10]  (.D(\input_filter[3][1] [10]), .CK(n_55_9), 
      .Q(\buffer[3][3][1] [10]), .QN());
   DFF_X1 \buffer_reg[3][3][1][9]  (.D(\input_filter[3][1] [9]), .CK(n_55_9), 
      .Q(\buffer[3][3][1] [9]), .QN());
   DFF_X1 \buffer_reg[3][3][1][8]  (.D(\input_filter[3][1] [8]), .CK(n_55_9), 
      .Q(\buffer[3][3][1] [8]), .QN());
   DFF_X1 \buffer_reg[3][3][1][7]  (.D(\input_filter[3][1] [7]), .CK(n_55_9), 
      .Q(\buffer[3][3][1] [7]), .QN());
   DFF_X1 \buffer_reg[3][3][1][6]  (.D(\input_filter[3][1] [6]), .CK(n_55_9), 
      .Q(\buffer[3][3][1] [6]), .QN());
   DFF_X1 \buffer_reg[3][3][1][5]  (.D(\input_filter[3][1] [5]), .CK(n_55_9), 
      .Q(\buffer[3][3][1] [5]), .QN());
   DFF_X1 \buffer_reg[3][3][1][4]  (.D(\input_filter[3][1] [4]), .CK(n_55_9), 
      .Q(\buffer[3][3][1] [4]), .QN());
   DFF_X1 \buffer_reg[3][3][1][3]  (.D(\input_filter[3][1] [3]), .CK(n_55_9), 
      .Q(\buffer[3][3][1] [3]), .QN());
   DFF_X1 \buffer_reg[3][3][1][2]  (.D(\input_filter[3][1] [2]), .CK(n_55_9), 
      .Q(\buffer[3][3][1] [2]), .QN());
   DFF_X1 \buffer_reg[3][3][1][1]  (.D(\input_filter[3][1] [1]), .CK(n_55_9), 
      .Q(\buffer[3][3][1] [1]), .QN());
   DFF_X1 \buffer_reg[3][3][1][0]  (.D(\input_filter[3][1] [0]), .CK(n_55_9), 
      .Q(\buffer[3][3][1] [0]), .QN());
   DFF_X1 \buffer_reg[2][3][1][15]  (.D(\input_filter[3][1] [15]), .CK(n_55_10), 
      .Q(\buffer[2][3][1] [15]), .QN());
   DFF_X1 \buffer_reg[2][3][1][14]  (.D(\input_filter[3][1] [14]), .CK(n_55_10), 
      .Q(\buffer[2][3][1] [14]), .QN());
   DFF_X1 \buffer_reg[2][3][1][13]  (.D(\input_filter[3][1] [13]), .CK(n_55_10), 
      .Q(\buffer[2][3][1] [13]), .QN());
   DFF_X1 \buffer_reg[2][3][1][12]  (.D(\input_filter[3][1] [12]), .CK(n_55_10), 
      .Q(\buffer[2][3][1] [12]), .QN());
   DFF_X1 \buffer_reg[2][3][1][11]  (.D(\input_filter[3][1] [11]), .CK(n_55_10), 
      .Q(\buffer[2][3][1] [11]), .QN());
   DFF_X1 \buffer_reg[2][3][1][10]  (.D(\input_filter[3][1] [10]), .CK(n_55_10), 
      .Q(\buffer[2][3][1] [10]), .QN());
   DFF_X1 \buffer_reg[2][3][1][9]  (.D(\input_filter[3][1] [9]), .CK(n_55_10), 
      .Q(\buffer[2][3][1] [9]), .QN());
   DFF_X1 \buffer_reg[2][3][1][8]  (.D(\input_filter[3][1] [8]), .CK(n_55_10), 
      .Q(\buffer[2][3][1] [8]), .QN());
   DFF_X1 \buffer_reg[2][3][1][7]  (.D(\input_filter[3][1] [7]), .CK(n_55_10), 
      .Q(\buffer[2][3][1] [7]), .QN());
   DFF_X1 \buffer_reg[2][3][1][6]  (.D(\input_filter[3][1] [6]), .CK(n_55_10), 
      .Q(\buffer[2][3][1] [6]), .QN());
   DFF_X1 \buffer_reg[2][3][1][5]  (.D(\input_filter[3][1] [5]), .CK(n_55_10), 
      .Q(\buffer[2][3][1] [5]), .QN());
   DFF_X1 \buffer_reg[2][3][1][4]  (.D(\input_filter[3][1] [4]), .CK(n_55_10), 
      .Q(\buffer[2][3][1] [4]), .QN());
   DFF_X1 \buffer_reg[2][3][1][3]  (.D(\input_filter[3][1] [3]), .CK(n_55_10), 
      .Q(\buffer[2][3][1] [3]), .QN());
   DFF_X1 \buffer_reg[2][3][1][2]  (.D(\input_filter[3][1] [2]), .CK(n_55_10), 
      .Q(\buffer[2][3][1] [2]), .QN());
   DFF_X1 \buffer_reg[2][3][1][1]  (.D(\input_filter[3][1] [1]), .CK(n_55_10), 
      .Q(\buffer[2][3][1] [1]), .QN());
   DFF_X1 \buffer_reg[2][3][1][0]  (.D(\input_filter[3][1] [0]), .CK(n_55_10), 
      .Q(\buffer[2][3][1] [0]), .QN());
   DFF_X1 \buffer_reg[1][3][1][15]  (.D(\input_filter[3][1] [15]), .CK(n_55_11), 
      .Q(\buffer[1][3][1] [15]), .QN());
   DFF_X1 \buffer_reg[1][3][1][14]  (.D(\input_filter[3][1] [14]), .CK(n_55_11), 
      .Q(\buffer[1][3][1] [14]), .QN());
   DFF_X1 \buffer_reg[1][3][1][13]  (.D(\input_filter[3][1] [13]), .CK(n_55_11), 
      .Q(\buffer[1][3][1] [13]), .QN());
   DFF_X1 \buffer_reg[1][3][1][12]  (.D(\input_filter[3][1] [12]), .CK(n_55_11), 
      .Q(\buffer[1][3][1] [12]), .QN());
   DFF_X1 \buffer_reg[1][3][1][11]  (.D(\input_filter[3][1] [11]), .CK(n_55_11), 
      .Q(\buffer[1][3][1] [11]), .QN());
   DFF_X1 \buffer_reg[1][3][1][10]  (.D(\input_filter[3][1] [10]), .CK(n_55_11), 
      .Q(\buffer[1][3][1] [10]), .QN());
   DFF_X1 \buffer_reg[1][3][1][9]  (.D(\input_filter[3][1] [9]), .CK(n_55_11), 
      .Q(\buffer[1][3][1] [9]), .QN());
   DFF_X1 \buffer_reg[1][3][1][8]  (.D(\input_filter[3][1] [8]), .CK(n_55_11), 
      .Q(\buffer[1][3][1] [8]), .QN());
   DFF_X1 \buffer_reg[1][3][1][7]  (.D(\input_filter[3][1] [7]), .CK(n_55_11), 
      .Q(\buffer[1][3][1] [7]), .QN());
   DFF_X1 \buffer_reg[1][3][1][6]  (.D(\input_filter[3][1] [6]), .CK(n_55_11), 
      .Q(\buffer[1][3][1] [6]), .QN());
   DFF_X1 \buffer_reg[1][3][1][5]  (.D(\input_filter[3][1] [5]), .CK(n_55_11), 
      .Q(\buffer[1][3][1] [5]), .QN());
   DFF_X1 \buffer_reg[1][3][1][4]  (.D(\input_filter[3][1] [4]), .CK(n_55_11), 
      .Q(\buffer[1][3][1] [4]), .QN());
   DFF_X1 \buffer_reg[1][3][1][3]  (.D(\input_filter[3][1] [3]), .CK(n_55_11), 
      .Q(\buffer[1][3][1] [3]), .QN());
   DFF_X1 \buffer_reg[1][3][1][2]  (.D(\input_filter[3][1] [2]), .CK(n_55_11), 
      .Q(\buffer[1][3][1] [2]), .QN());
   DFF_X1 \buffer_reg[1][3][1][1]  (.D(\input_filter[3][1] [1]), .CK(n_55_11), 
      .Q(\buffer[1][3][1] [1]), .QN());
   DFF_X1 \buffer_reg[1][3][1][0]  (.D(\input_filter[3][1] [0]), .CK(n_55_11), 
      .Q(\buffer[1][3][1] [0]), .QN());
   DFF_X1 \buffer_reg[0][3][1][15]  (.D(\input_filter[3][1] [15]), .CK(n_55_12), 
      .Q(\buffer[0][3][1] [15]), .QN());
   DFF_X1 \buffer_reg[0][3][1][14]  (.D(\input_filter[3][1] [14]), .CK(n_55_12), 
      .Q(\buffer[0][3][1] [14]), .QN());
   DFF_X1 \buffer_reg[0][3][1][13]  (.D(\input_filter[3][1] [13]), .CK(n_55_12), 
      .Q(\buffer[0][3][1] [13]), .QN());
   DFF_X1 \buffer_reg[0][3][1][12]  (.D(\input_filter[3][1] [12]), .CK(n_55_12), 
      .Q(\buffer[0][3][1] [12]), .QN());
   DFF_X1 \buffer_reg[0][3][1][11]  (.D(\input_filter[3][1] [11]), .CK(n_55_12), 
      .Q(\buffer[0][3][1] [11]), .QN());
   DFF_X1 \buffer_reg[0][3][1][10]  (.D(\input_filter[3][1] [10]), .CK(n_55_12), 
      .Q(\buffer[0][3][1] [10]), .QN());
   DFF_X1 \buffer_reg[0][3][1][9]  (.D(\input_filter[3][1] [9]), .CK(n_55_12), 
      .Q(\buffer[0][3][1] [9]), .QN());
   DFF_X1 \buffer_reg[0][3][1][8]  (.D(\input_filter[3][1] [8]), .CK(n_55_12), 
      .Q(\buffer[0][3][1] [8]), .QN());
   DFF_X1 \buffer_reg[0][3][1][7]  (.D(\input_filter[3][1] [7]), .CK(n_55_12), 
      .Q(\buffer[0][3][1] [7]), .QN());
   DFF_X1 \buffer_reg[0][3][1][6]  (.D(\input_filter[3][1] [6]), .CK(n_55_12), 
      .Q(\buffer[0][3][1] [6]), .QN());
   DFF_X1 \buffer_reg[0][3][1][5]  (.D(\input_filter[3][1] [5]), .CK(n_55_12), 
      .Q(\buffer[0][3][1] [5]), .QN());
   DFF_X1 \buffer_reg[0][3][1][4]  (.D(\input_filter[3][1] [4]), .CK(n_55_12), 
      .Q(\buffer[0][3][1] [4]), .QN());
   DFF_X1 \buffer_reg[0][3][1][3]  (.D(\input_filter[3][1] [3]), .CK(n_55_12), 
      .Q(\buffer[0][3][1] [3]), .QN());
   DFF_X1 \buffer_reg[0][3][1][2]  (.D(\input_filter[3][1] [2]), .CK(n_55_12), 
      .Q(\buffer[0][3][1] [2]), .QN());
   DFF_X1 \buffer_reg[0][3][1][1]  (.D(\input_filter[3][1] [1]), .CK(n_55_12), 
      .Q(\buffer[0][3][1] [1]), .QN());
   DFF_X1 \buffer_reg[0][3][1][0]  (.D(\input_filter[3][1] [0]), .CK(n_55_12), 
      .Q(\buffer[0][3][1] [0]), .QN());
   DFF_X1 \buffer_reg[15][3][0][15]  (.D(\input_filter[3][0] [15]), .CK(n_55_13), 
      .Q(\buffer[15][3][0] [15]), .QN());
   DFF_X1 \buffer_reg[15][3][0][14]  (.D(\input_filter[3][0] [14]), .CK(n_55_13), 
      .Q(\buffer[15][3][0] [14]), .QN());
   DFF_X1 \buffer_reg[15][3][0][13]  (.D(\input_filter[3][0] [13]), .CK(n_55_13), 
      .Q(\buffer[15][3][0] [13]), .QN());
   DFF_X1 \buffer_reg[15][3][0][12]  (.D(\input_filter[3][0] [12]), .CK(n_55_13), 
      .Q(\buffer[15][3][0] [12]), .QN());
   DFF_X1 \buffer_reg[15][3][0][11]  (.D(\input_filter[3][0] [11]), .CK(n_55_13), 
      .Q(\buffer[15][3][0] [11]), .QN());
   DFF_X1 \buffer_reg[15][3][0][10]  (.D(\input_filter[3][0] [10]), .CK(n_55_13), 
      .Q(\buffer[15][3][0] [10]), .QN());
   DFF_X1 \buffer_reg[15][3][0][9]  (.D(\input_filter[3][0] [9]), .CK(n_55_13), 
      .Q(\buffer[15][3][0] [9]), .QN());
   DFF_X1 \buffer_reg[15][3][0][8]  (.D(\input_filter[3][0] [8]), .CK(n_55_13), 
      .Q(\buffer[15][3][0] [8]), .QN());
   DFF_X1 \buffer_reg[15][3][0][7]  (.D(\input_filter[3][0] [7]), .CK(n_55_13), 
      .Q(\buffer[15][3][0] [7]), .QN());
   DFF_X1 \buffer_reg[15][3][0][6]  (.D(\input_filter[3][0] [6]), .CK(n_55_13), 
      .Q(\buffer[15][3][0] [6]), .QN());
   DFF_X1 \buffer_reg[15][3][0][5]  (.D(\input_filter[3][0] [5]), .CK(n_55_13), 
      .Q(\buffer[15][3][0] [5]), .QN());
   DFF_X1 \buffer_reg[15][3][0][4]  (.D(\input_filter[3][0] [4]), .CK(n_55_13), 
      .Q(\buffer[15][3][0] [4]), .QN());
   DFF_X1 \buffer_reg[15][3][0][3]  (.D(\input_filter[3][0] [3]), .CK(n_55_13), 
      .Q(\buffer[15][3][0] [3]), .QN());
   DFF_X1 \buffer_reg[15][3][0][2]  (.D(\input_filter[3][0] [2]), .CK(n_55_13), 
      .Q(\buffer[15][3][0] [2]), .QN());
   DFF_X1 \buffer_reg[15][3][0][1]  (.D(\input_filter[3][0] [1]), .CK(n_55_13), 
      .Q(\buffer[15][3][0] [1]), .QN());
   DFF_X1 \buffer_reg[15][3][0][0]  (.D(\input_filter[3][0] [0]), .CK(n_55_13), 
      .Q(\buffer[15][3][0] [0]), .QN());
   DFF_X1 \buffer_reg[14][3][0][15]  (.D(\input_filter[3][0] [15]), .CK(n_55_14), 
      .Q(\buffer[14][3][0] [15]), .QN());
   DFF_X1 \buffer_reg[14][3][0][14]  (.D(\input_filter[3][0] [14]), .CK(n_55_14), 
      .Q(\buffer[14][3][0] [14]), .QN());
   DFF_X1 \buffer_reg[14][3][0][13]  (.D(\input_filter[3][0] [13]), .CK(n_55_14), 
      .Q(\buffer[14][3][0] [13]), .QN());
   DFF_X1 \buffer_reg[14][3][0][12]  (.D(\input_filter[3][0] [12]), .CK(n_55_14), 
      .Q(\buffer[14][3][0] [12]), .QN());
   DFF_X1 \buffer_reg[14][3][0][11]  (.D(\input_filter[3][0] [11]), .CK(n_55_14), 
      .Q(\buffer[14][3][0] [11]), .QN());
   DFF_X1 \buffer_reg[14][3][0][10]  (.D(\input_filter[3][0] [10]), .CK(n_55_14), 
      .Q(\buffer[14][3][0] [10]), .QN());
   DFF_X1 \buffer_reg[14][3][0][9]  (.D(\input_filter[3][0] [9]), .CK(n_55_14), 
      .Q(\buffer[14][3][0] [9]), .QN());
   DFF_X1 \buffer_reg[14][3][0][8]  (.D(\input_filter[3][0] [8]), .CK(n_55_14), 
      .Q(\buffer[14][3][0] [8]), .QN());
   DFF_X1 \buffer_reg[14][3][0][7]  (.D(\input_filter[3][0] [7]), .CK(n_55_14), 
      .Q(\buffer[14][3][0] [7]), .QN());
   DFF_X1 \buffer_reg[14][3][0][6]  (.D(\input_filter[3][0] [6]), .CK(n_55_14), 
      .Q(\buffer[14][3][0] [6]), .QN());
   DFF_X1 \buffer_reg[14][3][0][5]  (.D(\input_filter[3][0] [5]), .CK(n_55_14), 
      .Q(\buffer[14][3][0] [5]), .QN());
   DFF_X1 \buffer_reg[14][3][0][4]  (.D(\input_filter[3][0] [4]), .CK(n_55_14), 
      .Q(\buffer[14][3][0] [4]), .QN());
   DFF_X1 \buffer_reg[14][3][0][3]  (.D(\input_filter[3][0] [3]), .CK(n_55_14), 
      .Q(\buffer[14][3][0] [3]), .QN());
   DFF_X1 \buffer_reg[14][3][0][2]  (.D(\input_filter[3][0] [2]), .CK(n_55_14), 
      .Q(\buffer[14][3][0] [2]), .QN());
   DFF_X1 \buffer_reg[14][3][0][1]  (.D(\input_filter[3][0] [1]), .CK(n_55_14), 
      .Q(\buffer[14][3][0] [1]), .QN());
   DFF_X1 \buffer_reg[14][3][0][0]  (.D(\input_filter[3][0] [0]), .CK(n_55_14), 
      .Q(\buffer[14][3][0] [0]), .QN());
   DFF_X1 \buffer_reg[13][3][0][15]  (.D(\input_filter[3][0] [15]), .CK(n_55_15), 
      .Q(\buffer[13][3][0] [15]), .QN());
   DFF_X1 \buffer_reg[13][3][0][14]  (.D(\input_filter[3][0] [14]), .CK(n_55_15), 
      .Q(\buffer[13][3][0] [14]), .QN());
   DFF_X1 \buffer_reg[13][3][0][13]  (.D(\input_filter[3][0] [13]), .CK(n_55_15), 
      .Q(\buffer[13][3][0] [13]), .QN());
   DFF_X1 \buffer_reg[13][3][0][12]  (.D(\input_filter[3][0] [12]), .CK(n_55_15), 
      .Q(\buffer[13][3][0] [12]), .QN());
   DFF_X1 \buffer_reg[13][3][0][11]  (.D(\input_filter[3][0] [11]), .CK(n_55_15), 
      .Q(\buffer[13][3][0] [11]), .QN());
   DFF_X1 \buffer_reg[13][3][0][10]  (.D(\input_filter[3][0] [10]), .CK(n_55_15), 
      .Q(\buffer[13][3][0] [10]), .QN());
   DFF_X1 \buffer_reg[13][3][0][9]  (.D(\input_filter[3][0] [9]), .CK(n_55_15), 
      .Q(\buffer[13][3][0] [9]), .QN());
   DFF_X1 \buffer_reg[13][3][0][8]  (.D(\input_filter[3][0] [8]), .CK(n_55_15), 
      .Q(\buffer[13][3][0] [8]), .QN());
   DFF_X1 \buffer_reg[13][3][0][7]  (.D(\input_filter[3][0] [7]), .CK(n_55_15), 
      .Q(\buffer[13][3][0] [7]), .QN());
   DFF_X1 \buffer_reg[13][3][0][6]  (.D(\input_filter[3][0] [6]), .CK(n_55_15), 
      .Q(\buffer[13][3][0] [6]), .QN());
   DFF_X1 \buffer_reg[13][3][0][5]  (.D(\input_filter[3][0] [5]), .CK(n_55_15), 
      .Q(\buffer[13][3][0] [5]), .QN());
   DFF_X1 \buffer_reg[13][3][0][4]  (.D(\input_filter[3][0] [4]), .CK(n_55_15), 
      .Q(\buffer[13][3][0] [4]), .QN());
   DFF_X1 \buffer_reg[13][3][0][3]  (.D(\input_filter[3][0] [3]), .CK(n_55_15), 
      .Q(\buffer[13][3][0] [3]), .QN());
   DFF_X1 \buffer_reg[13][3][0][2]  (.D(\input_filter[3][0] [2]), .CK(n_55_15), 
      .Q(\buffer[13][3][0] [2]), .QN());
   DFF_X1 \buffer_reg[13][3][0][1]  (.D(\input_filter[3][0] [1]), .CK(n_55_15), 
      .Q(\buffer[13][3][0] [1]), .QN());
   DFF_X1 \buffer_reg[13][3][0][0]  (.D(\input_filter[3][0] [0]), .CK(n_55_15), 
      .Q(\buffer[13][3][0] [0]), .QN());
   DFF_X1 \buffer_reg[12][3][0][15]  (.D(\input_filter[3][0] [15]), .CK(n_55_0), 
      .Q(\buffer[12][3][0] [15]), .QN());
   DFF_X1 \buffer_reg[12][3][0][14]  (.D(\input_filter[3][0] [14]), .CK(n_55_0), 
      .Q(\buffer[12][3][0] [14]), .QN());
   DFF_X1 \buffer_reg[12][3][0][13]  (.D(\input_filter[3][0] [13]), .CK(n_55_0), 
      .Q(\buffer[12][3][0] [13]), .QN());
   DFF_X1 \buffer_reg[12][3][0][12]  (.D(\input_filter[3][0] [12]), .CK(n_55_0), 
      .Q(\buffer[12][3][0] [12]), .QN());
   DFF_X1 \buffer_reg[12][3][0][11]  (.D(\input_filter[3][0] [11]), .CK(n_55_0), 
      .Q(\buffer[12][3][0] [11]), .QN());
   DFF_X1 \buffer_reg[12][3][0][10]  (.D(\input_filter[3][0] [10]), .CK(n_55_0), 
      .Q(\buffer[12][3][0] [10]), .QN());
   DFF_X1 \buffer_reg[12][3][0][9]  (.D(\input_filter[3][0] [9]), .CK(n_55_0), 
      .Q(\buffer[12][3][0] [9]), .QN());
   DFF_X1 \buffer_reg[12][3][0][8]  (.D(\input_filter[3][0] [8]), .CK(n_55_0), 
      .Q(\buffer[12][3][0] [8]), .QN());
   DFF_X1 \buffer_reg[12][3][0][7]  (.D(\input_filter[3][0] [7]), .CK(n_55_0), 
      .Q(\buffer[12][3][0] [7]), .QN());
   DFF_X1 \buffer_reg[12][3][0][6]  (.D(\input_filter[3][0] [6]), .CK(n_55_0), 
      .Q(\buffer[12][3][0] [6]), .QN());
   DFF_X1 \buffer_reg[12][3][0][5]  (.D(\input_filter[3][0] [5]), .CK(n_55_0), 
      .Q(\buffer[12][3][0] [5]), .QN());
   DFF_X1 \buffer_reg[12][3][0][4]  (.D(\input_filter[3][0] [4]), .CK(n_55_0), 
      .Q(\buffer[12][3][0] [4]), .QN());
   DFF_X1 \buffer_reg[12][3][0][3]  (.D(\input_filter[3][0] [3]), .CK(n_55_0), 
      .Q(\buffer[12][3][0] [3]), .QN());
   DFF_X1 \buffer_reg[12][3][0][2]  (.D(\input_filter[3][0] [2]), .CK(n_55_0), 
      .Q(\buffer[12][3][0] [2]), .QN());
   DFF_X1 \buffer_reg[12][3][0][1]  (.D(\input_filter[3][0] [1]), .CK(n_55_0), 
      .Q(\buffer[12][3][0] [1]), .QN());
   DFF_X1 \buffer_reg[12][3][0][0]  (.D(\input_filter[3][0] [0]), .CK(n_55_0), 
      .Q(\buffer[12][3][0] [0]), .QN());
   DFF_X1 \buffer_reg[11][3][0][15]  (.D(\input_filter[3][0] [15]), .CK(n_55_1), 
      .Q(\buffer[11][3][0] [15]), .QN());
   DFF_X1 \buffer_reg[11][3][0][14]  (.D(\input_filter[3][0] [14]), .CK(n_55_1), 
      .Q(\buffer[11][3][0] [14]), .QN());
   DFF_X1 \buffer_reg[11][3][0][13]  (.D(\input_filter[3][0] [13]), .CK(n_55_1), 
      .Q(\buffer[11][3][0] [13]), .QN());
   DFF_X1 \buffer_reg[11][3][0][12]  (.D(\input_filter[3][0] [12]), .CK(n_55_1), 
      .Q(\buffer[11][3][0] [12]), .QN());
   DFF_X1 \buffer_reg[11][3][0][11]  (.D(\input_filter[3][0] [11]), .CK(n_55_1), 
      .Q(\buffer[11][3][0] [11]), .QN());
   DFF_X1 \buffer_reg[11][3][0][10]  (.D(\input_filter[3][0] [10]), .CK(n_55_1), 
      .Q(\buffer[11][3][0] [10]), .QN());
   DFF_X1 \buffer_reg[11][3][0][9]  (.D(\input_filter[3][0] [9]), .CK(n_55_1), 
      .Q(\buffer[11][3][0] [9]), .QN());
   DFF_X1 \buffer_reg[11][3][0][8]  (.D(\input_filter[3][0] [8]), .CK(n_55_1), 
      .Q(\buffer[11][3][0] [8]), .QN());
   DFF_X1 \buffer_reg[11][3][0][7]  (.D(\input_filter[3][0] [7]), .CK(n_55_1), 
      .Q(\buffer[11][3][0] [7]), .QN());
   DFF_X1 \buffer_reg[11][3][0][6]  (.D(\input_filter[3][0] [6]), .CK(n_55_1), 
      .Q(\buffer[11][3][0] [6]), .QN());
   DFF_X1 \buffer_reg[11][3][0][5]  (.D(\input_filter[3][0] [5]), .CK(n_55_1), 
      .Q(\buffer[11][3][0] [5]), .QN());
   DFF_X1 \buffer_reg[11][3][0][4]  (.D(\input_filter[3][0] [4]), .CK(n_55_1), 
      .Q(\buffer[11][3][0] [4]), .QN());
   DFF_X1 \buffer_reg[11][3][0][3]  (.D(\input_filter[3][0] [3]), .CK(n_55_1), 
      .Q(\buffer[11][3][0] [3]), .QN());
   DFF_X1 \buffer_reg[11][3][0][2]  (.D(\input_filter[3][0] [2]), .CK(n_55_1), 
      .Q(\buffer[11][3][0] [2]), .QN());
   DFF_X1 \buffer_reg[11][3][0][1]  (.D(\input_filter[3][0] [1]), .CK(n_55_1), 
      .Q(\buffer[11][3][0] [1]), .QN());
   DFF_X1 \buffer_reg[11][3][0][0]  (.D(\input_filter[3][0] [0]), .CK(n_55_1), 
      .Q(\buffer[11][3][0] [0]), .QN());
   DFF_X1 \buffer_reg[10][3][0][15]  (.D(\input_filter[3][0] [15]), .CK(n_55_2), 
      .Q(\buffer[10][3][0] [15]), .QN());
   DFF_X1 \buffer_reg[10][3][0][14]  (.D(\input_filter[3][0] [14]), .CK(n_55_2), 
      .Q(\buffer[10][3][0] [14]), .QN());
   DFF_X1 \buffer_reg[10][3][0][13]  (.D(\input_filter[3][0] [13]), .CK(n_55_2), 
      .Q(\buffer[10][3][0] [13]), .QN());
   DFF_X1 \buffer_reg[10][3][0][12]  (.D(\input_filter[3][0] [12]), .CK(n_55_2), 
      .Q(\buffer[10][3][0] [12]), .QN());
   DFF_X1 \buffer_reg[10][3][0][11]  (.D(\input_filter[3][0] [11]), .CK(n_55_2), 
      .Q(\buffer[10][3][0] [11]), .QN());
   DFF_X1 \buffer_reg[10][3][0][10]  (.D(\input_filter[3][0] [10]), .CK(n_55_2), 
      .Q(\buffer[10][3][0] [10]), .QN());
   DFF_X1 \buffer_reg[10][3][0][9]  (.D(\input_filter[3][0] [9]), .CK(n_55_2), 
      .Q(\buffer[10][3][0] [9]), .QN());
   DFF_X1 \buffer_reg[10][3][0][8]  (.D(\input_filter[3][0] [8]), .CK(n_55_2), 
      .Q(\buffer[10][3][0] [8]), .QN());
   DFF_X1 \buffer_reg[10][3][0][7]  (.D(\input_filter[3][0] [7]), .CK(n_55_2), 
      .Q(\buffer[10][3][0] [7]), .QN());
   DFF_X1 \buffer_reg[10][3][0][6]  (.D(\input_filter[3][0] [6]), .CK(n_55_2), 
      .Q(\buffer[10][3][0] [6]), .QN());
   DFF_X1 \buffer_reg[10][3][0][5]  (.D(\input_filter[3][0] [5]), .CK(n_55_2), 
      .Q(\buffer[10][3][0] [5]), .QN());
   DFF_X1 \buffer_reg[10][3][0][4]  (.D(\input_filter[3][0] [4]), .CK(n_55_2), 
      .Q(\buffer[10][3][0] [4]), .QN());
   DFF_X1 \buffer_reg[10][3][0][3]  (.D(\input_filter[3][0] [3]), .CK(n_55_2), 
      .Q(\buffer[10][3][0] [3]), .QN());
   DFF_X1 \buffer_reg[10][3][0][2]  (.D(\input_filter[3][0] [2]), .CK(n_55_2), 
      .Q(\buffer[10][3][0] [2]), .QN());
   DFF_X1 \buffer_reg[10][3][0][1]  (.D(\input_filter[3][0] [1]), .CK(n_55_2), 
      .Q(\buffer[10][3][0] [1]), .QN());
   DFF_X1 \buffer_reg[10][3][0][0]  (.D(\input_filter[3][0] [0]), .CK(n_55_2), 
      .Q(\buffer[10][3][0] [0]), .QN());
   DFF_X1 \buffer_reg[9][3][0][15]  (.D(\input_filter[3][0] [15]), .CK(n_55_3), 
      .Q(\buffer[9][3][0] [15]), .QN());
   DFF_X1 \buffer_reg[9][3][0][14]  (.D(\input_filter[3][0] [14]), .CK(n_55_3), 
      .Q(\buffer[9][3][0] [14]), .QN());
   DFF_X1 \buffer_reg[9][3][0][13]  (.D(\input_filter[3][0] [13]), .CK(n_55_3), 
      .Q(\buffer[9][3][0] [13]), .QN());
   DFF_X1 \buffer_reg[9][3][0][12]  (.D(\input_filter[3][0] [12]), .CK(n_55_3), 
      .Q(\buffer[9][3][0] [12]), .QN());
   DFF_X1 \buffer_reg[9][3][0][11]  (.D(\input_filter[3][0] [11]), .CK(n_55_3), 
      .Q(\buffer[9][3][0] [11]), .QN());
   DFF_X1 \buffer_reg[9][3][0][10]  (.D(\input_filter[3][0] [10]), .CK(n_55_3), 
      .Q(\buffer[9][3][0] [10]), .QN());
   DFF_X1 \buffer_reg[9][3][0][9]  (.D(\input_filter[3][0] [9]), .CK(n_55_3), 
      .Q(\buffer[9][3][0] [9]), .QN());
   DFF_X1 \buffer_reg[9][3][0][8]  (.D(\input_filter[3][0] [8]), .CK(n_55_3), 
      .Q(\buffer[9][3][0] [8]), .QN());
   DFF_X1 \buffer_reg[9][3][0][7]  (.D(\input_filter[3][0] [7]), .CK(n_55_3), 
      .Q(\buffer[9][3][0] [7]), .QN());
   DFF_X1 \buffer_reg[9][3][0][6]  (.D(\input_filter[3][0] [6]), .CK(n_55_3), 
      .Q(\buffer[9][3][0] [6]), .QN());
   DFF_X1 \buffer_reg[9][3][0][5]  (.D(\input_filter[3][0] [5]), .CK(n_55_3), 
      .Q(\buffer[9][3][0] [5]), .QN());
   DFF_X1 \buffer_reg[9][3][0][4]  (.D(\input_filter[3][0] [4]), .CK(n_55_3), 
      .Q(\buffer[9][3][0] [4]), .QN());
   DFF_X1 \buffer_reg[9][3][0][3]  (.D(\input_filter[3][0] [3]), .CK(n_55_3), 
      .Q(\buffer[9][3][0] [3]), .QN());
   DFF_X1 \buffer_reg[9][3][0][2]  (.D(\input_filter[3][0] [2]), .CK(n_55_3), 
      .Q(\buffer[9][3][0] [2]), .QN());
   DFF_X1 \buffer_reg[9][3][0][1]  (.D(\input_filter[3][0] [1]), .CK(n_55_3), 
      .Q(\buffer[9][3][0] [1]), .QN());
   DFF_X1 \buffer_reg[9][3][0][0]  (.D(\input_filter[3][0] [0]), .CK(n_55_3), 
      .Q(\buffer[9][3][0] [0]), .QN());
   DFF_X1 \buffer_reg[8][3][0][15]  (.D(\input_filter[3][0] [15]), .CK(n_55_4), 
      .Q(\buffer[8][3][0] [15]), .QN());
   DFF_X1 \buffer_reg[8][3][0][14]  (.D(\input_filter[3][0] [14]), .CK(n_55_4), 
      .Q(\buffer[8][3][0] [14]), .QN());
   DFF_X1 \buffer_reg[8][3][0][13]  (.D(\input_filter[3][0] [13]), .CK(n_55_4), 
      .Q(\buffer[8][3][0] [13]), .QN());
   DFF_X1 \buffer_reg[8][3][0][12]  (.D(\input_filter[3][0] [12]), .CK(n_55_4), 
      .Q(\buffer[8][3][0] [12]), .QN());
   DFF_X1 \buffer_reg[8][3][0][11]  (.D(\input_filter[3][0] [11]), .CK(n_55_4), 
      .Q(\buffer[8][3][0] [11]), .QN());
   DFF_X1 \buffer_reg[8][3][0][10]  (.D(\input_filter[3][0] [10]), .CK(n_55_4), 
      .Q(\buffer[8][3][0] [10]), .QN());
   DFF_X1 \buffer_reg[8][3][0][9]  (.D(\input_filter[3][0] [9]), .CK(n_55_4), 
      .Q(\buffer[8][3][0] [9]), .QN());
   DFF_X1 \buffer_reg[8][3][0][8]  (.D(\input_filter[3][0] [8]), .CK(n_55_4), 
      .Q(\buffer[8][3][0] [8]), .QN());
   DFF_X1 \buffer_reg[8][3][0][7]  (.D(\input_filter[3][0] [7]), .CK(n_55_4), 
      .Q(\buffer[8][3][0] [7]), .QN());
   DFF_X1 \buffer_reg[8][3][0][6]  (.D(\input_filter[3][0] [6]), .CK(n_55_4), 
      .Q(\buffer[8][3][0] [6]), .QN());
   DFF_X1 \buffer_reg[8][3][0][5]  (.D(\input_filter[3][0] [5]), .CK(n_55_4), 
      .Q(\buffer[8][3][0] [5]), .QN());
   DFF_X1 \buffer_reg[8][3][0][4]  (.D(\input_filter[3][0] [4]), .CK(n_55_4), 
      .Q(\buffer[8][3][0] [4]), .QN());
   DFF_X1 \buffer_reg[8][3][0][3]  (.D(\input_filter[3][0] [3]), .CK(n_55_4), 
      .Q(\buffer[8][3][0] [3]), .QN());
   DFF_X1 \buffer_reg[8][3][0][2]  (.D(\input_filter[3][0] [2]), .CK(n_55_4), 
      .Q(\buffer[8][3][0] [2]), .QN());
   DFF_X1 \buffer_reg[8][3][0][1]  (.D(\input_filter[3][0] [1]), .CK(n_55_4), 
      .Q(\buffer[8][3][0] [1]), .QN());
   DFF_X1 \buffer_reg[8][3][0][0]  (.D(\input_filter[3][0] [0]), .CK(n_55_4), 
      .Q(\buffer[8][3][0] [0]), .QN());
   DFF_X1 \buffer_reg[7][3][0][15]  (.D(\input_filter[3][0] [15]), .CK(n_55_5), 
      .Q(\buffer[7][3][0] [15]), .QN());
   DFF_X1 \buffer_reg[7][3][0][14]  (.D(\input_filter[3][0] [14]), .CK(n_55_5), 
      .Q(\buffer[7][3][0] [14]), .QN());
   DFF_X1 \buffer_reg[7][3][0][13]  (.D(\input_filter[3][0] [13]), .CK(n_55_5), 
      .Q(\buffer[7][3][0] [13]), .QN());
   DFF_X1 \buffer_reg[7][3][0][12]  (.D(\input_filter[3][0] [12]), .CK(n_55_5), 
      .Q(\buffer[7][3][0] [12]), .QN());
   DFF_X1 \buffer_reg[7][3][0][11]  (.D(\input_filter[3][0] [11]), .CK(n_55_5), 
      .Q(\buffer[7][3][0] [11]), .QN());
   DFF_X1 \buffer_reg[7][3][0][10]  (.D(\input_filter[3][0] [10]), .CK(n_55_5), 
      .Q(\buffer[7][3][0] [10]), .QN());
   DFF_X1 \buffer_reg[7][3][0][9]  (.D(\input_filter[3][0] [9]), .CK(n_55_5), 
      .Q(\buffer[7][3][0] [9]), .QN());
   DFF_X1 \buffer_reg[7][3][0][8]  (.D(\input_filter[3][0] [8]), .CK(n_55_5), 
      .Q(\buffer[7][3][0] [8]), .QN());
   DFF_X1 \buffer_reg[7][3][0][7]  (.D(\input_filter[3][0] [7]), .CK(n_55_5), 
      .Q(\buffer[7][3][0] [7]), .QN());
   DFF_X1 \buffer_reg[7][3][0][6]  (.D(\input_filter[3][0] [6]), .CK(n_55_5), 
      .Q(\buffer[7][3][0] [6]), .QN());
   DFF_X1 \buffer_reg[7][3][0][5]  (.D(\input_filter[3][0] [5]), .CK(n_55_5), 
      .Q(\buffer[7][3][0] [5]), .QN());
   DFF_X1 \buffer_reg[7][3][0][4]  (.D(\input_filter[3][0] [4]), .CK(n_55_5), 
      .Q(\buffer[7][3][0] [4]), .QN());
   DFF_X1 \buffer_reg[7][3][0][3]  (.D(\input_filter[3][0] [3]), .CK(n_55_5), 
      .Q(\buffer[7][3][0] [3]), .QN());
   DFF_X1 \buffer_reg[7][3][0][2]  (.D(\input_filter[3][0] [2]), .CK(n_55_5), 
      .Q(\buffer[7][3][0] [2]), .QN());
   DFF_X1 \buffer_reg[7][3][0][1]  (.D(\input_filter[3][0] [1]), .CK(n_55_5), 
      .Q(\buffer[7][3][0] [1]), .QN());
   DFF_X1 \buffer_reg[7][3][0][0]  (.D(\input_filter[3][0] [0]), .CK(n_55_5), 
      .Q(\buffer[7][3][0] [0]), .QN());
   DFF_X1 \buffer_reg[6][3][0][15]  (.D(\input_filter[3][0] [15]), .CK(n_55_6), 
      .Q(\buffer[6][3][0] [15]), .QN());
   DFF_X1 \buffer_reg[6][3][0][14]  (.D(\input_filter[3][0] [14]), .CK(n_55_6), 
      .Q(\buffer[6][3][0] [14]), .QN());
   DFF_X1 \buffer_reg[6][3][0][13]  (.D(\input_filter[3][0] [13]), .CK(n_55_6), 
      .Q(\buffer[6][3][0] [13]), .QN());
   DFF_X1 \buffer_reg[6][3][0][12]  (.D(\input_filter[3][0] [12]), .CK(n_55_6), 
      .Q(\buffer[6][3][0] [12]), .QN());
   DFF_X1 \buffer_reg[6][3][0][11]  (.D(\input_filter[3][0] [11]), .CK(n_55_6), 
      .Q(\buffer[6][3][0] [11]), .QN());
   DFF_X1 \buffer_reg[6][3][0][10]  (.D(\input_filter[3][0] [10]), .CK(n_55_6), 
      .Q(\buffer[6][3][0] [10]), .QN());
   DFF_X1 \buffer_reg[6][3][0][9]  (.D(\input_filter[3][0] [9]), .CK(n_55_6), 
      .Q(\buffer[6][3][0] [9]), .QN());
   DFF_X1 \buffer_reg[6][3][0][8]  (.D(\input_filter[3][0] [8]), .CK(n_55_6), 
      .Q(\buffer[6][3][0] [8]), .QN());
   DFF_X1 \buffer_reg[6][3][0][7]  (.D(\input_filter[3][0] [7]), .CK(n_55_6), 
      .Q(\buffer[6][3][0] [7]), .QN());
   DFF_X1 \buffer_reg[6][3][0][6]  (.D(\input_filter[3][0] [6]), .CK(n_55_6), 
      .Q(\buffer[6][3][0] [6]), .QN());
   DFF_X1 \buffer_reg[6][3][0][5]  (.D(\input_filter[3][0] [5]), .CK(n_55_6), 
      .Q(\buffer[6][3][0] [5]), .QN());
   DFF_X1 \buffer_reg[6][3][0][4]  (.D(\input_filter[3][0] [4]), .CK(n_55_6), 
      .Q(\buffer[6][3][0] [4]), .QN());
   DFF_X1 \buffer_reg[6][3][0][3]  (.D(\input_filter[3][0] [3]), .CK(n_55_6), 
      .Q(\buffer[6][3][0] [3]), .QN());
   DFF_X1 \buffer_reg[6][3][0][2]  (.D(\input_filter[3][0] [2]), .CK(n_55_6), 
      .Q(\buffer[6][3][0] [2]), .QN());
   DFF_X1 \buffer_reg[6][3][0][1]  (.D(\input_filter[3][0] [1]), .CK(n_55_6), 
      .Q(\buffer[6][3][0] [1]), .QN());
   DFF_X1 \buffer_reg[6][3][0][0]  (.D(\input_filter[3][0] [0]), .CK(n_55_6), 
      .Q(\buffer[6][3][0] [0]), .QN());
   DFF_X1 \buffer_reg[5][3][0][15]  (.D(\input_filter[3][0] [15]), .CK(n_55_7), 
      .Q(\buffer[5][3][0] [15]), .QN());
   DFF_X1 \buffer_reg[5][3][0][14]  (.D(\input_filter[3][0] [14]), .CK(n_55_7), 
      .Q(\buffer[5][3][0] [14]), .QN());
   DFF_X1 \buffer_reg[5][3][0][13]  (.D(\input_filter[3][0] [13]), .CK(n_55_7), 
      .Q(\buffer[5][3][0] [13]), .QN());
   DFF_X1 \buffer_reg[5][3][0][12]  (.D(\input_filter[3][0] [12]), .CK(n_55_7), 
      .Q(\buffer[5][3][0] [12]), .QN());
   DFF_X1 \buffer_reg[5][3][0][11]  (.D(\input_filter[3][0] [11]), .CK(n_55_7), 
      .Q(\buffer[5][3][0] [11]), .QN());
   DFF_X1 \buffer_reg[5][3][0][10]  (.D(\input_filter[3][0] [10]), .CK(n_55_7), 
      .Q(\buffer[5][3][0] [10]), .QN());
   DFF_X1 \buffer_reg[5][3][0][9]  (.D(\input_filter[3][0] [9]), .CK(n_55_7), 
      .Q(\buffer[5][3][0] [9]), .QN());
   DFF_X1 \buffer_reg[5][3][0][8]  (.D(\input_filter[3][0] [8]), .CK(n_55_7), 
      .Q(\buffer[5][3][0] [8]), .QN());
   DFF_X1 \buffer_reg[5][3][0][7]  (.D(\input_filter[3][0] [7]), .CK(n_55_7), 
      .Q(\buffer[5][3][0] [7]), .QN());
   DFF_X1 \buffer_reg[5][3][0][6]  (.D(\input_filter[3][0] [6]), .CK(n_55_7), 
      .Q(\buffer[5][3][0] [6]), .QN());
   DFF_X1 \buffer_reg[5][3][0][5]  (.D(\input_filter[3][0] [5]), .CK(n_55_7), 
      .Q(\buffer[5][3][0] [5]), .QN());
   DFF_X1 \buffer_reg[5][3][0][4]  (.D(\input_filter[3][0] [4]), .CK(n_55_7), 
      .Q(\buffer[5][3][0] [4]), .QN());
   DFF_X1 \buffer_reg[5][3][0][3]  (.D(\input_filter[3][0] [3]), .CK(n_55_7), 
      .Q(\buffer[5][3][0] [3]), .QN());
   DFF_X1 \buffer_reg[5][3][0][2]  (.D(\input_filter[3][0] [2]), .CK(n_55_7), 
      .Q(\buffer[5][3][0] [2]), .QN());
   DFF_X1 \buffer_reg[5][3][0][1]  (.D(\input_filter[3][0] [1]), .CK(n_55_7), 
      .Q(\buffer[5][3][0] [1]), .QN());
   DFF_X1 \buffer_reg[5][3][0][0]  (.D(\input_filter[3][0] [0]), .CK(n_55_7), 
      .Q(\buffer[5][3][0] [0]), .QN());
   DFF_X1 \buffer_reg[4][3][0][15]  (.D(\input_filter[3][0] [15]), .CK(n_55_8), 
      .Q(\buffer[4][3][0] [15]), .QN());
   DFF_X1 \buffer_reg[4][3][0][14]  (.D(\input_filter[3][0] [14]), .CK(n_55_8), 
      .Q(\buffer[4][3][0] [14]), .QN());
   DFF_X1 \buffer_reg[4][3][0][13]  (.D(\input_filter[3][0] [13]), .CK(n_55_8), 
      .Q(\buffer[4][3][0] [13]), .QN());
   DFF_X1 \buffer_reg[4][3][0][12]  (.D(\input_filter[3][0] [12]), .CK(n_55_8), 
      .Q(\buffer[4][3][0] [12]), .QN());
   DFF_X1 \buffer_reg[4][3][0][11]  (.D(\input_filter[3][0] [11]), .CK(n_55_8), 
      .Q(\buffer[4][3][0] [11]), .QN());
   DFF_X1 \buffer_reg[4][3][0][10]  (.D(\input_filter[3][0] [10]), .CK(n_55_8), 
      .Q(\buffer[4][3][0] [10]), .QN());
   DFF_X1 \buffer_reg[4][3][0][9]  (.D(\input_filter[3][0] [9]), .CK(n_55_8), 
      .Q(\buffer[4][3][0] [9]), .QN());
   DFF_X1 \buffer_reg[4][3][0][8]  (.D(\input_filter[3][0] [8]), .CK(n_55_8), 
      .Q(\buffer[4][3][0] [8]), .QN());
   DFF_X1 \buffer_reg[4][3][0][7]  (.D(\input_filter[3][0] [7]), .CK(n_55_8), 
      .Q(\buffer[4][3][0] [7]), .QN());
   DFF_X1 \buffer_reg[4][3][0][6]  (.D(\input_filter[3][0] [6]), .CK(n_55_8), 
      .Q(\buffer[4][3][0] [6]), .QN());
   DFF_X1 \buffer_reg[4][3][0][5]  (.D(\input_filter[3][0] [5]), .CK(n_55_8), 
      .Q(\buffer[4][3][0] [5]), .QN());
   DFF_X1 \buffer_reg[4][3][0][4]  (.D(\input_filter[3][0] [4]), .CK(n_55_8), 
      .Q(\buffer[4][3][0] [4]), .QN());
   DFF_X1 \buffer_reg[4][3][0][3]  (.D(\input_filter[3][0] [3]), .CK(n_55_8), 
      .Q(\buffer[4][3][0] [3]), .QN());
   DFF_X1 \buffer_reg[4][3][0][2]  (.D(\input_filter[3][0] [2]), .CK(n_55_8), 
      .Q(\buffer[4][3][0] [2]), .QN());
   DFF_X1 \buffer_reg[4][3][0][1]  (.D(\input_filter[3][0] [1]), .CK(n_55_8), 
      .Q(\buffer[4][3][0] [1]), .QN());
   DFF_X1 \buffer_reg[4][3][0][0]  (.D(\input_filter[3][0] [0]), .CK(n_55_8), 
      .Q(\buffer[4][3][0] [0]), .QN());
   DFF_X1 \buffer_reg[3][3][0][15]  (.D(\input_filter[3][0] [15]), .CK(n_55_9), 
      .Q(\buffer[3][3][0] [15]), .QN());
   DFF_X1 \buffer_reg[3][3][0][14]  (.D(\input_filter[3][0] [14]), .CK(n_55_9), 
      .Q(\buffer[3][3][0] [14]), .QN());
   DFF_X1 \buffer_reg[3][3][0][13]  (.D(\input_filter[3][0] [13]), .CK(n_55_9), 
      .Q(\buffer[3][3][0] [13]), .QN());
   DFF_X1 \buffer_reg[3][3][0][12]  (.D(\input_filter[3][0] [12]), .CK(n_55_9), 
      .Q(\buffer[3][3][0] [12]), .QN());
   DFF_X1 \buffer_reg[3][3][0][11]  (.D(\input_filter[3][0] [11]), .CK(n_55_9), 
      .Q(\buffer[3][3][0] [11]), .QN());
   DFF_X1 \buffer_reg[3][3][0][10]  (.D(\input_filter[3][0] [10]), .CK(n_55_9), 
      .Q(\buffer[3][3][0] [10]), .QN());
   DFF_X1 \buffer_reg[3][3][0][9]  (.D(\input_filter[3][0] [9]), .CK(n_55_9), 
      .Q(\buffer[3][3][0] [9]), .QN());
   DFF_X1 \buffer_reg[3][3][0][8]  (.D(\input_filter[3][0] [8]), .CK(n_55_9), 
      .Q(\buffer[3][3][0] [8]), .QN());
   DFF_X1 \buffer_reg[3][3][0][7]  (.D(\input_filter[3][0] [7]), .CK(n_55_9), 
      .Q(\buffer[3][3][0] [7]), .QN());
   DFF_X1 \buffer_reg[3][3][0][6]  (.D(\input_filter[3][0] [6]), .CK(n_55_9), 
      .Q(\buffer[3][3][0] [6]), .QN());
   DFF_X1 \buffer_reg[3][3][0][5]  (.D(\input_filter[3][0] [5]), .CK(n_55_9), 
      .Q(\buffer[3][3][0] [5]), .QN());
   DFF_X1 \buffer_reg[3][3][0][4]  (.D(\input_filter[3][0] [4]), .CK(n_55_9), 
      .Q(\buffer[3][3][0] [4]), .QN());
   DFF_X1 \buffer_reg[3][3][0][3]  (.D(\input_filter[3][0] [3]), .CK(n_55_9), 
      .Q(\buffer[3][3][0] [3]), .QN());
   DFF_X1 \buffer_reg[3][3][0][2]  (.D(\input_filter[3][0] [2]), .CK(n_55_9), 
      .Q(\buffer[3][3][0] [2]), .QN());
   DFF_X1 \buffer_reg[3][3][0][1]  (.D(\input_filter[3][0] [1]), .CK(n_55_9), 
      .Q(\buffer[3][3][0] [1]), .QN());
   DFF_X1 \buffer_reg[3][3][0][0]  (.D(\input_filter[3][0] [0]), .CK(n_55_9), 
      .Q(\buffer[3][3][0] [0]), .QN());
   DFF_X1 \buffer_reg[2][3][0][15]  (.D(\input_filter[3][0] [15]), .CK(n_55_10), 
      .Q(\buffer[2][3][0] [15]), .QN());
   DFF_X1 \buffer_reg[2][3][0][14]  (.D(\input_filter[3][0] [14]), .CK(n_55_10), 
      .Q(\buffer[2][3][0] [14]), .QN());
   DFF_X1 \buffer_reg[2][3][0][13]  (.D(\input_filter[3][0] [13]), .CK(n_55_10), 
      .Q(\buffer[2][3][0] [13]), .QN());
   DFF_X1 \buffer_reg[2][3][0][12]  (.D(\input_filter[3][0] [12]), .CK(n_55_10), 
      .Q(\buffer[2][3][0] [12]), .QN());
   DFF_X1 \buffer_reg[2][3][0][11]  (.D(\input_filter[3][0] [11]), .CK(n_55_10), 
      .Q(\buffer[2][3][0] [11]), .QN());
   DFF_X1 \buffer_reg[2][3][0][10]  (.D(\input_filter[3][0] [10]), .CK(n_55_10), 
      .Q(\buffer[2][3][0] [10]), .QN());
   DFF_X1 \buffer_reg[2][3][0][9]  (.D(\input_filter[3][0] [9]), .CK(n_55_10), 
      .Q(\buffer[2][3][0] [9]), .QN());
   DFF_X1 \buffer_reg[2][3][0][8]  (.D(\input_filter[3][0] [8]), .CK(n_55_10), 
      .Q(\buffer[2][3][0] [8]), .QN());
   DFF_X1 \buffer_reg[2][3][0][7]  (.D(\input_filter[3][0] [7]), .CK(n_55_10), 
      .Q(\buffer[2][3][0] [7]), .QN());
   DFF_X1 \buffer_reg[2][3][0][6]  (.D(\input_filter[3][0] [6]), .CK(n_55_10), 
      .Q(\buffer[2][3][0] [6]), .QN());
   DFF_X1 \buffer_reg[2][3][0][5]  (.D(\input_filter[3][0] [5]), .CK(n_55_10), 
      .Q(\buffer[2][3][0] [5]), .QN());
   DFF_X1 \buffer_reg[2][3][0][4]  (.D(\input_filter[3][0] [4]), .CK(n_55_10), 
      .Q(\buffer[2][3][0] [4]), .QN());
   DFF_X1 \buffer_reg[2][3][0][3]  (.D(\input_filter[3][0] [3]), .CK(n_55_10), 
      .Q(\buffer[2][3][0] [3]), .QN());
   DFF_X1 \buffer_reg[2][3][0][2]  (.D(\input_filter[3][0] [2]), .CK(n_55_10), 
      .Q(\buffer[2][3][0] [2]), .QN());
   DFF_X1 \buffer_reg[2][3][0][1]  (.D(\input_filter[3][0] [1]), .CK(n_55_10), 
      .Q(\buffer[2][3][0] [1]), .QN());
   DFF_X1 \buffer_reg[2][3][0][0]  (.D(\input_filter[3][0] [0]), .CK(n_55_10), 
      .Q(\buffer[2][3][0] [0]), .QN());
   DFF_X1 \buffer_reg[1][3][0][15]  (.D(\input_filter[3][0] [15]), .CK(n_55_11), 
      .Q(\buffer[1][3][0] [15]), .QN());
   DFF_X1 \buffer_reg[1][3][0][14]  (.D(\input_filter[3][0] [14]), .CK(n_55_11), 
      .Q(\buffer[1][3][0] [14]), .QN());
   DFF_X1 \buffer_reg[1][3][0][13]  (.D(\input_filter[3][0] [13]), .CK(n_55_11), 
      .Q(\buffer[1][3][0] [13]), .QN());
   DFF_X1 \buffer_reg[1][3][0][12]  (.D(\input_filter[3][0] [12]), .CK(n_55_11), 
      .Q(\buffer[1][3][0] [12]), .QN());
   DFF_X1 \buffer_reg[1][3][0][11]  (.D(\input_filter[3][0] [11]), .CK(n_55_11), 
      .Q(\buffer[1][3][0] [11]), .QN());
   DFF_X1 \buffer_reg[1][3][0][10]  (.D(\input_filter[3][0] [10]), .CK(n_55_11), 
      .Q(\buffer[1][3][0] [10]), .QN());
   DFF_X1 \buffer_reg[1][3][0][9]  (.D(\input_filter[3][0] [9]), .CK(n_55_11), 
      .Q(\buffer[1][3][0] [9]), .QN());
   DFF_X1 \buffer_reg[1][3][0][8]  (.D(\input_filter[3][0] [8]), .CK(n_55_11), 
      .Q(\buffer[1][3][0] [8]), .QN());
   DFF_X1 \buffer_reg[1][3][0][7]  (.D(\input_filter[3][0] [7]), .CK(n_55_11), 
      .Q(\buffer[1][3][0] [7]), .QN());
   DFF_X1 \buffer_reg[1][3][0][6]  (.D(\input_filter[3][0] [6]), .CK(n_55_11), 
      .Q(\buffer[1][3][0] [6]), .QN());
   DFF_X1 \buffer_reg[1][3][0][5]  (.D(\input_filter[3][0] [5]), .CK(n_55_11), 
      .Q(\buffer[1][3][0] [5]), .QN());
   DFF_X1 \buffer_reg[1][3][0][4]  (.D(\input_filter[3][0] [4]), .CK(n_55_11), 
      .Q(\buffer[1][3][0] [4]), .QN());
   DFF_X1 \buffer_reg[1][3][0][3]  (.D(\input_filter[3][0] [3]), .CK(n_55_11), 
      .Q(\buffer[1][3][0] [3]), .QN());
   DFF_X1 \buffer_reg[1][3][0][2]  (.D(\input_filter[3][0] [2]), .CK(n_55_11), 
      .Q(\buffer[1][3][0] [2]), .QN());
   DFF_X1 \buffer_reg[1][3][0][1]  (.D(\input_filter[3][0] [1]), .CK(n_55_11), 
      .Q(\buffer[1][3][0] [1]), .QN());
   DFF_X1 \buffer_reg[1][3][0][0]  (.D(\input_filter[3][0] [0]), .CK(n_55_11), 
      .Q(\buffer[1][3][0] [0]), .QN());
   DFF_X1 \buffer_reg[0][3][0][15]  (.D(\input_filter[3][0] [15]), .CK(n_55_12), 
      .Q(\buffer[0][3][0] [15]), .QN());
   DFF_X1 \buffer_reg[0][3][0][14]  (.D(\input_filter[3][0] [14]), .CK(n_55_12), 
      .Q(\buffer[0][3][0] [14]), .QN());
   DFF_X1 \buffer_reg[0][3][0][13]  (.D(\input_filter[3][0] [13]), .CK(n_55_12), 
      .Q(\buffer[0][3][0] [13]), .QN());
   DFF_X1 \buffer_reg[0][3][0][12]  (.D(\input_filter[3][0] [12]), .CK(n_55_12), 
      .Q(\buffer[0][3][0] [12]), .QN());
   DFF_X1 \buffer_reg[0][3][0][11]  (.D(\input_filter[3][0] [11]), .CK(n_55_12), 
      .Q(\buffer[0][3][0] [11]), .QN());
   DFF_X1 \buffer_reg[0][3][0][10]  (.D(\input_filter[3][0] [10]), .CK(n_55_12), 
      .Q(\buffer[0][3][0] [10]), .QN());
   DFF_X1 \buffer_reg[0][3][0][9]  (.D(\input_filter[3][0] [9]), .CK(n_55_12), 
      .Q(\buffer[0][3][0] [9]), .QN());
   DFF_X1 \buffer_reg[0][3][0][8]  (.D(\input_filter[3][0] [8]), .CK(n_55_12), 
      .Q(\buffer[0][3][0] [8]), .QN());
   DFF_X1 \buffer_reg[0][3][0][7]  (.D(\input_filter[3][0] [7]), .CK(n_55_12), 
      .Q(\buffer[0][3][0] [7]), .QN());
   DFF_X1 \buffer_reg[0][3][0][6]  (.D(\input_filter[3][0] [6]), .CK(n_55_12), 
      .Q(\buffer[0][3][0] [6]), .QN());
   DFF_X1 \buffer_reg[0][3][0][5]  (.D(\input_filter[3][0] [5]), .CK(n_55_12), 
      .Q(\buffer[0][3][0] [5]), .QN());
   DFF_X1 \buffer_reg[0][3][0][4]  (.D(\input_filter[3][0] [4]), .CK(n_55_12), 
      .Q(\buffer[0][3][0] [4]), .QN());
   DFF_X1 \buffer_reg[0][3][0][3]  (.D(\input_filter[3][0] [3]), .CK(n_55_12), 
      .Q(\buffer[0][3][0] [3]), .QN());
   DFF_X1 \buffer_reg[0][3][0][2]  (.D(\input_filter[3][0] [2]), .CK(n_55_12), 
      .Q(\buffer[0][3][0] [2]), .QN());
   DFF_X1 \buffer_reg[0][3][0][1]  (.D(\input_filter[3][0] [1]), .CK(n_55_12), 
      .Q(\buffer[0][3][0] [1]), .QN());
   DFF_X1 \buffer_reg[0][3][0][0]  (.D(\input_filter[3][0] [0]), .CK(n_55_12), 
      .Q(\buffer[0][3][0] [0]), .QN());
   DFF_X1 \buffer_reg[15][2][4][15]  (.D(\input_filter[2][4] [15]), .CK(n_55_13), 
      .Q(\buffer[15][2][4] [15]), .QN());
   DFF_X1 \buffer_reg[15][2][4][14]  (.D(\input_filter[2][4] [14]), .CK(n_55_13), 
      .Q(\buffer[15][2][4] [14]), .QN());
   DFF_X1 \buffer_reg[15][2][4][13]  (.D(\input_filter[2][4] [13]), .CK(n_55_13), 
      .Q(\buffer[15][2][4] [13]), .QN());
   DFF_X1 \buffer_reg[15][2][4][12]  (.D(\input_filter[2][4] [12]), .CK(n_55_13), 
      .Q(\buffer[15][2][4] [12]), .QN());
   DFF_X1 \buffer_reg[15][2][4][11]  (.D(\input_filter[2][4] [11]), .CK(n_55_13), 
      .Q(\buffer[15][2][4] [11]), .QN());
   DFF_X1 \buffer_reg[15][2][4][10]  (.D(\input_filter[2][4] [10]), .CK(n_55_13), 
      .Q(\buffer[15][2][4] [10]), .QN());
   DFF_X1 \buffer_reg[15][2][4][9]  (.D(\input_filter[2][4] [9]), .CK(n_55_13), 
      .Q(\buffer[15][2][4] [9]), .QN());
   DFF_X1 \buffer_reg[15][2][4][8]  (.D(\input_filter[2][4] [8]), .CK(n_55_13), 
      .Q(\buffer[15][2][4] [8]), .QN());
   DFF_X1 \buffer_reg[15][2][4][7]  (.D(\input_filter[2][4] [7]), .CK(n_55_13), 
      .Q(\buffer[15][2][4] [7]), .QN());
   DFF_X1 \buffer_reg[15][2][4][6]  (.D(\input_filter[2][4] [6]), .CK(n_55_13), 
      .Q(\buffer[15][2][4] [6]), .QN());
   DFF_X1 \buffer_reg[15][2][4][5]  (.D(\input_filter[2][4] [5]), .CK(n_55_13), 
      .Q(\buffer[15][2][4] [5]), .QN());
   DFF_X1 \buffer_reg[15][2][4][4]  (.D(\input_filter[2][4] [4]), .CK(n_55_13), 
      .Q(\buffer[15][2][4] [4]), .QN());
   DFF_X1 \buffer_reg[15][2][4][3]  (.D(\input_filter[2][4] [3]), .CK(n_55_13), 
      .Q(\buffer[15][2][4] [3]), .QN());
   DFF_X1 \buffer_reg[15][2][4][2]  (.D(\input_filter[2][4] [2]), .CK(n_55_13), 
      .Q(\buffer[15][2][4] [2]), .QN());
   DFF_X1 \buffer_reg[15][2][4][1]  (.D(\input_filter[2][4] [1]), .CK(n_55_13), 
      .Q(\buffer[15][2][4] [1]), .QN());
   DFF_X1 \buffer_reg[15][2][4][0]  (.D(\input_filter[2][4] [0]), .CK(n_55_13), 
      .Q(\buffer[15][2][4] [0]), .QN());
   DFF_X1 \buffer_reg[14][2][4][15]  (.D(\input_filter[2][4] [15]), .CK(n_55_14), 
      .Q(\buffer[14][2][4] [15]), .QN());
   DFF_X1 \buffer_reg[14][2][4][14]  (.D(\input_filter[2][4] [14]), .CK(n_55_14), 
      .Q(\buffer[14][2][4] [14]), .QN());
   DFF_X1 \buffer_reg[14][2][4][13]  (.D(\input_filter[2][4] [13]), .CK(n_55_14), 
      .Q(\buffer[14][2][4] [13]), .QN());
   DFF_X1 \buffer_reg[14][2][4][12]  (.D(\input_filter[2][4] [12]), .CK(n_55_14), 
      .Q(\buffer[14][2][4] [12]), .QN());
   DFF_X1 \buffer_reg[14][2][4][11]  (.D(\input_filter[2][4] [11]), .CK(n_55_14), 
      .Q(\buffer[14][2][4] [11]), .QN());
   DFF_X1 \buffer_reg[14][2][4][10]  (.D(\input_filter[2][4] [10]), .CK(n_55_14), 
      .Q(\buffer[14][2][4] [10]), .QN());
   DFF_X1 \buffer_reg[14][2][4][9]  (.D(\input_filter[2][4] [9]), .CK(n_55_14), 
      .Q(\buffer[14][2][4] [9]), .QN());
   DFF_X1 \buffer_reg[14][2][4][8]  (.D(\input_filter[2][4] [8]), .CK(n_55_14), 
      .Q(\buffer[14][2][4] [8]), .QN());
   DFF_X1 \buffer_reg[14][2][4][7]  (.D(\input_filter[2][4] [7]), .CK(n_55_14), 
      .Q(\buffer[14][2][4] [7]), .QN());
   DFF_X1 \buffer_reg[14][2][4][6]  (.D(\input_filter[2][4] [6]), .CK(n_55_14), 
      .Q(\buffer[14][2][4] [6]), .QN());
   DFF_X1 \buffer_reg[14][2][4][5]  (.D(\input_filter[2][4] [5]), .CK(n_55_14), 
      .Q(\buffer[14][2][4] [5]), .QN());
   DFF_X1 \buffer_reg[14][2][4][4]  (.D(\input_filter[2][4] [4]), .CK(n_55_14), 
      .Q(\buffer[14][2][4] [4]), .QN());
   DFF_X1 \buffer_reg[14][2][4][3]  (.D(\input_filter[2][4] [3]), .CK(n_55_14), 
      .Q(\buffer[14][2][4] [3]), .QN());
   DFF_X1 \buffer_reg[14][2][4][2]  (.D(\input_filter[2][4] [2]), .CK(n_55_14), 
      .Q(\buffer[14][2][4] [2]), .QN());
   DFF_X1 \buffer_reg[14][2][4][1]  (.D(\input_filter[2][4] [1]), .CK(n_55_14), 
      .Q(\buffer[14][2][4] [1]), .QN());
   DFF_X1 \buffer_reg[14][2][4][0]  (.D(\input_filter[2][4] [0]), .CK(n_55_14), 
      .Q(\buffer[14][2][4] [0]), .QN());
   DFF_X1 \buffer_reg[13][2][4][15]  (.D(\input_filter[2][4] [15]), .CK(n_55_15), 
      .Q(\buffer[13][2][4] [15]), .QN());
   DFF_X1 \buffer_reg[13][2][4][14]  (.D(\input_filter[2][4] [14]), .CK(n_55_15), 
      .Q(\buffer[13][2][4] [14]), .QN());
   DFF_X1 \buffer_reg[13][2][4][13]  (.D(\input_filter[2][4] [13]), .CK(n_55_15), 
      .Q(\buffer[13][2][4] [13]), .QN());
   DFF_X1 \buffer_reg[13][2][4][12]  (.D(\input_filter[2][4] [12]), .CK(n_55_15), 
      .Q(\buffer[13][2][4] [12]), .QN());
   DFF_X1 \buffer_reg[13][2][4][11]  (.D(\input_filter[2][4] [11]), .CK(n_55_15), 
      .Q(\buffer[13][2][4] [11]), .QN());
   DFF_X1 \buffer_reg[13][2][4][10]  (.D(\input_filter[2][4] [10]), .CK(n_55_15), 
      .Q(\buffer[13][2][4] [10]), .QN());
   DFF_X1 \buffer_reg[13][2][4][9]  (.D(\input_filter[2][4] [9]), .CK(n_55_15), 
      .Q(\buffer[13][2][4] [9]), .QN());
   DFF_X1 \buffer_reg[13][2][4][8]  (.D(\input_filter[2][4] [8]), .CK(n_55_15), 
      .Q(\buffer[13][2][4] [8]), .QN());
   DFF_X1 \buffer_reg[13][2][4][7]  (.D(\input_filter[2][4] [7]), .CK(n_55_15), 
      .Q(\buffer[13][2][4] [7]), .QN());
   DFF_X1 \buffer_reg[13][2][4][6]  (.D(\input_filter[2][4] [6]), .CK(n_55_15), 
      .Q(\buffer[13][2][4] [6]), .QN());
   DFF_X1 \buffer_reg[13][2][4][5]  (.D(\input_filter[2][4] [5]), .CK(n_55_15), 
      .Q(\buffer[13][2][4] [5]), .QN());
   DFF_X1 \buffer_reg[13][2][4][4]  (.D(\input_filter[2][4] [4]), .CK(n_55_15), 
      .Q(\buffer[13][2][4] [4]), .QN());
   DFF_X1 \buffer_reg[13][2][4][3]  (.D(\input_filter[2][4] [3]), .CK(n_55_15), 
      .Q(\buffer[13][2][4] [3]), .QN());
   DFF_X1 \buffer_reg[13][2][4][2]  (.D(\input_filter[2][4] [2]), .CK(n_55_15), 
      .Q(\buffer[13][2][4] [2]), .QN());
   DFF_X1 \buffer_reg[13][2][4][1]  (.D(\input_filter[2][4] [1]), .CK(n_55_15), 
      .Q(\buffer[13][2][4] [1]), .QN());
   DFF_X1 \buffer_reg[13][2][4][0]  (.D(\input_filter[2][4] [0]), .CK(n_55_15), 
      .Q(\buffer[13][2][4] [0]), .QN());
   DFF_X1 \buffer_reg[12][2][4][15]  (.D(\input_filter[2][4] [15]), .CK(n_55_0), 
      .Q(\buffer[12][2][4] [15]), .QN());
   DFF_X1 \buffer_reg[12][2][4][14]  (.D(\input_filter[2][4] [14]), .CK(n_55_0), 
      .Q(\buffer[12][2][4] [14]), .QN());
   DFF_X1 \buffer_reg[12][2][4][13]  (.D(\input_filter[2][4] [13]), .CK(n_55_0), 
      .Q(\buffer[12][2][4] [13]), .QN());
   DFF_X1 \buffer_reg[12][2][4][12]  (.D(\input_filter[2][4] [12]), .CK(n_55_0), 
      .Q(\buffer[12][2][4] [12]), .QN());
   DFF_X1 \buffer_reg[12][2][4][11]  (.D(\input_filter[2][4] [11]), .CK(n_55_0), 
      .Q(\buffer[12][2][4] [11]), .QN());
   DFF_X1 \buffer_reg[12][2][4][10]  (.D(\input_filter[2][4] [10]), .CK(n_55_0), 
      .Q(\buffer[12][2][4] [10]), .QN());
   DFF_X1 \buffer_reg[12][2][4][9]  (.D(\input_filter[2][4] [9]), .CK(n_55_0), 
      .Q(\buffer[12][2][4] [9]), .QN());
   DFF_X1 \buffer_reg[12][2][4][8]  (.D(\input_filter[2][4] [8]), .CK(n_55_0), 
      .Q(\buffer[12][2][4] [8]), .QN());
   DFF_X1 \buffer_reg[12][2][4][7]  (.D(\input_filter[2][4] [7]), .CK(n_55_0), 
      .Q(\buffer[12][2][4] [7]), .QN());
   DFF_X1 \buffer_reg[12][2][4][6]  (.D(\input_filter[2][4] [6]), .CK(n_55_0), 
      .Q(\buffer[12][2][4] [6]), .QN());
   DFF_X1 \buffer_reg[12][2][4][5]  (.D(\input_filter[2][4] [5]), .CK(n_55_0), 
      .Q(\buffer[12][2][4] [5]), .QN());
   DFF_X1 \buffer_reg[12][2][4][4]  (.D(\input_filter[2][4] [4]), .CK(n_55_0), 
      .Q(\buffer[12][2][4] [4]), .QN());
   DFF_X1 \buffer_reg[12][2][4][3]  (.D(\input_filter[2][4] [3]), .CK(n_55_0), 
      .Q(\buffer[12][2][4] [3]), .QN());
   DFF_X1 \buffer_reg[12][2][4][2]  (.D(\input_filter[2][4] [2]), .CK(n_55_0), 
      .Q(\buffer[12][2][4] [2]), .QN());
   DFF_X1 \buffer_reg[12][2][4][1]  (.D(\input_filter[2][4] [1]), .CK(n_55_0), 
      .Q(\buffer[12][2][4] [1]), .QN());
   DFF_X1 \buffer_reg[12][2][4][0]  (.D(\input_filter[2][4] [0]), .CK(n_55_0), 
      .Q(\buffer[12][2][4] [0]), .QN());
   DFF_X1 \buffer_reg[11][2][4][15]  (.D(\input_filter[2][4] [15]), .CK(n_55_1), 
      .Q(\buffer[11][2][4] [15]), .QN());
   DFF_X1 \buffer_reg[11][2][4][14]  (.D(\input_filter[2][4] [14]), .CK(n_55_1), 
      .Q(\buffer[11][2][4] [14]), .QN());
   DFF_X1 \buffer_reg[11][2][4][13]  (.D(\input_filter[2][4] [13]), .CK(n_55_1), 
      .Q(\buffer[11][2][4] [13]), .QN());
   DFF_X1 \buffer_reg[11][2][4][12]  (.D(\input_filter[2][4] [12]), .CK(n_55_1), 
      .Q(\buffer[11][2][4] [12]), .QN());
   DFF_X1 \buffer_reg[11][2][4][11]  (.D(\input_filter[2][4] [11]), .CK(n_55_1), 
      .Q(\buffer[11][2][4] [11]), .QN());
   DFF_X1 \buffer_reg[11][2][4][10]  (.D(\input_filter[2][4] [10]), .CK(n_55_1), 
      .Q(\buffer[11][2][4] [10]), .QN());
   DFF_X1 \buffer_reg[11][2][4][9]  (.D(\input_filter[2][4] [9]), .CK(n_55_1), 
      .Q(\buffer[11][2][4] [9]), .QN());
   DFF_X1 \buffer_reg[11][2][4][8]  (.D(\input_filter[2][4] [8]), .CK(n_55_1), 
      .Q(\buffer[11][2][4] [8]), .QN());
   DFF_X1 \buffer_reg[11][2][4][7]  (.D(\input_filter[2][4] [7]), .CK(n_55_1), 
      .Q(\buffer[11][2][4] [7]), .QN());
   DFF_X1 \buffer_reg[11][2][4][6]  (.D(\input_filter[2][4] [6]), .CK(n_55_1), 
      .Q(\buffer[11][2][4] [6]), .QN());
   DFF_X1 \buffer_reg[11][2][4][5]  (.D(\input_filter[2][4] [5]), .CK(n_55_1), 
      .Q(\buffer[11][2][4] [5]), .QN());
   DFF_X1 \buffer_reg[11][2][4][4]  (.D(\input_filter[2][4] [4]), .CK(n_55_1), 
      .Q(\buffer[11][2][4] [4]), .QN());
   DFF_X1 \buffer_reg[11][2][4][3]  (.D(\input_filter[2][4] [3]), .CK(n_55_1), 
      .Q(\buffer[11][2][4] [3]), .QN());
   DFF_X1 \buffer_reg[11][2][4][2]  (.D(\input_filter[2][4] [2]), .CK(n_55_1), 
      .Q(\buffer[11][2][4] [2]), .QN());
   DFF_X1 \buffer_reg[11][2][4][1]  (.D(\input_filter[2][4] [1]), .CK(n_55_1), 
      .Q(\buffer[11][2][4] [1]), .QN());
   DFF_X1 \buffer_reg[11][2][4][0]  (.D(\input_filter[2][4] [0]), .CK(n_55_1), 
      .Q(\buffer[11][2][4] [0]), .QN());
   DFF_X1 \buffer_reg[10][2][4][15]  (.D(\input_filter[2][4] [15]), .CK(n_55_2), 
      .Q(\buffer[10][2][4] [15]), .QN());
   DFF_X1 \buffer_reg[10][2][4][14]  (.D(\input_filter[2][4] [14]), .CK(n_55_2), 
      .Q(\buffer[10][2][4] [14]), .QN());
   DFF_X1 \buffer_reg[10][2][4][13]  (.D(\input_filter[2][4] [13]), .CK(n_55_2), 
      .Q(\buffer[10][2][4] [13]), .QN());
   DFF_X1 \buffer_reg[10][2][4][12]  (.D(\input_filter[2][4] [12]), .CK(n_55_2), 
      .Q(\buffer[10][2][4] [12]), .QN());
   DFF_X1 \buffer_reg[10][2][4][11]  (.D(\input_filter[2][4] [11]), .CK(n_55_2), 
      .Q(\buffer[10][2][4] [11]), .QN());
   DFF_X1 \buffer_reg[10][2][4][10]  (.D(\input_filter[2][4] [10]), .CK(n_55_2), 
      .Q(\buffer[10][2][4] [10]), .QN());
   DFF_X1 \buffer_reg[10][2][4][9]  (.D(\input_filter[2][4] [9]), .CK(n_55_2), 
      .Q(\buffer[10][2][4] [9]), .QN());
   DFF_X1 \buffer_reg[10][2][4][8]  (.D(\input_filter[2][4] [8]), .CK(n_55_2), 
      .Q(\buffer[10][2][4] [8]), .QN());
   DFF_X1 \buffer_reg[10][2][4][7]  (.D(\input_filter[2][4] [7]), .CK(n_55_2), 
      .Q(\buffer[10][2][4] [7]), .QN());
   DFF_X1 \buffer_reg[10][2][4][6]  (.D(\input_filter[2][4] [6]), .CK(n_55_2), 
      .Q(\buffer[10][2][4] [6]), .QN());
   DFF_X1 \buffer_reg[10][2][4][5]  (.D(\input_filter[2][4] [5]), .CK(n_55_2), 
      .Q(\buffer[10][2][4] [5]), .QN());
   DFF_X1 \buffer_reg[10][2][4][4]  (.D(\input_filter[2][4] [4]), .CK(n_55_2), 
      .Q(\buffer[10][2][4] [4]), .QN());
   DFF_X1 \buffer_reg[10][2][4][3]  (.D(\input_filter[2][4] [3]), .CK(n_55_2), 
      .Q(\buffer[10][2][4] [3]), .QN());
   DFF_X1 \buffer_reg[10][2][4][2]  (.D(\input_filter[2][4] [2]), .CK(n_55_2), 
      .Q(\buffer[10][2][4] [2]), .QN());
   DFF_X1 \buffer_reg[10][2][4][1]  (.D(\input_filter[2][4] [1]), .CK(n_55_2), 
      .Q(\buffer[10][2][4] [1]), .QN());
   DFF_X1 \buffer_reg[10][2][4][0]  (.D(\input_filter[2][4] [0]), .CK(n_55_2), 
      .Q(\buffer[10][2][4] [0]), .QN());
   DFF_X1 \buffer_reg[9][2][4][15]  (.D(\input_filter[2][4] [15]), .CK(n_55_3), 
      .Q(\buffer[9][2][4] [15]), .QN());
   DFF_X1 \buffer_reg[9][2][4][14]  (.D(\input_filter[2][4] [14]), .CK(n_55_3), 
      .Q(\buffer[9][2][4] [14]), .QN());
   DFF_X1 \buffer_reg[9][2][4][13]  (.D(\input_filter[2][4] [13]), .CK(n_55_3), 
      .Q(\buffer[9][2][4] [13]), .QN());
   DFF_X1 \buffer_reg[9][2][4][12]  (.D(\input_filter[2][4] [12]), .CK(n_55_3), 
      .Q(\buffer[9][2][4] [12]), .QN());
   DFF_X1 \buffer_reg[9][2][4][11]  (.D(\input_filter[2][4] [11]), .CK(n_55_3), 
      .Q(\buffer[9][2][4] [11]), .QN());
   DFF_X1 \buffer_reg[9][2][4][10]  (.D(\input_filter[2][4] [10]), .CK(n_55_3), 
      .Q(\buffer[9][2][4] [10]), .QN());
   DFF_X1 \buffer_reg[9][2][4][9]  (.D(\input_filter[2][4] [9]), .CK(n_55_3), 
      .Q(\buffer[9][2][4] [9]), .QN());
   DFF_X1 \buffer_reg[9][2][4][8]  (.D(\input_filter[2][4] [8]), .CK(n_55_3), 
      .Q(\buffer[9][2][4] [8]), .QN());
   DFF_X1 \buffer_reg[9][2][4][7]  (.D(\input_filter[2][4] [7]), .CK(n_55_3), 
      .Q(\buffer[9][2][4] [7]), .QN());
   DFF_X1 \buffer_reg[9][2][4][6]  (.D(\input_filter[2][4] [6]), .CK(n_55_3), 
      .Q(\buffer[9][2][4] [6]), .QN());
   DFF_X1 \buffer_reg[9][2][4][5]  (.D(\input_filter[2][4] [5]), .CK(n_55_3), 
      .Q(\buffer[9][2][4] [5]), .QN());
   DFF_X1 \buffer_reg[9][2][4][4]  (.D(\input_filter[2][4] [4]), .CK(n_55_3), 
      .Q(\buffer[9][2][4] [4]), .QN());
   DFF_X1 \buffer_reg[9][2][4][3]  (.D(\input_filter[2][4] [3]), .CK(n_55_3), 
      .Q(\buffer[9][2][4] [3]), .QN());
   DFF_X1 \buffer_reg[9][2][4][2]  (.D(\input_filter[2][4] [2]), .CK(n_55_3), 
      .Q(\buffer[9][2][4] [2]), .QN());
   DFF_X1 \buffer_reg[9][2][4][1]  (.D(\input_filter[2][4] [1]), .CK(n_55_3), 
      .Q(\buffer[9][2][4] [1]), .QN());
   DFF_X1 \buffer_reg[9][2][4][0]  (.D(\input_filter[2][4] [0]), .CK(n_55_3), 
      .Q(\buffer[9][2][4] [0]), .QN());
   DFF_X1 \buffer_reg[8][2][4][15]  (.D(\input_filter[2][4] [15]), .CK(n_55_4), 
      .Q(\buffer[8][2][4] [15]), .QN());
   DFF_X1 \buffer_reg[8][2][4][14]  (.D(\input_filter[2][4] [14]), .CK(n_55_4), 
      .Q(\buffer[8][2][4] [14]), .QN());
   DFF_X1 \buffer_reg[8][2][4][13]  (.D(\input_filter[2][4] [13]), .CK(n_55_4), 
      .Q(\buffer[8][2][4] [13]), .QN());
   DFF_X1 \buffer_reg[8][2][4][12]  (.D(\input_filter[2][4] [12]), .CK(n_55_4), 
      .Q(\buffer[8][2][4] [12]), .QN());
   DFF_X1 \buffer_reg[8][2][4][11]  (.D(\input_filter[2][4] [11]), .CK(n_55_4), 
      .Q(\buffer[8][2][4] [11]), .QN());
   DFF_X1 \buffer_reg[8][2][4][10]  (.D(\input_filter[2][4] [10]), .CK(n_55_4), 
      .Q(\buffer[8][2][4] [10]), .QN());
   DFF_X1 \buffer_reg[8][2][4][9]  (.D(\input_filter[2][4] [9]), .CK(n_55_4), 
      .Q(\buffer[8][2][4] [9]), .QN());
   DFF_X1 \buffer_reg[8][2][4][8]  (.D(\input_filter[2][4] [8]), .CK(n_55_4), 
      .Q(\buffer[8][2][4] [8]), .QN());
   DFF_X1 \buffer_reg[8][2][4][7]  (.D(\input_filter[2][4] [7]), .CK(n_55_4), 
      .Q(\buffer[8][2][4] [7]), .QN());
   DFF_X1 \buffer_reg[8][2][4][6]  (.D(\input_filter[2][4] [6]), .CK(n_55_4), 
      .Q(\buffer[8][2][4] [6]), .QN());
   DFF_X1 \buffer_reg[8][2][4][5]  (.D(\input_filter[2][4] [5]), .CK(n_55_4), 
      .Q(\buffer[8][2][4] [5]), .QN());
   DFF_X1 \buffer_reg[8][2][4][4]  (.D(\input_filter[2][4] [4]), .CK(n_55_4), 
      .Q(\buffer[8][2][4] [4]), .QN());
   DFF_X1 \buffer_reg[8][2][4][3]  (.D(\input_filter[2][4] [3]), .CK(n_55_4), 
      .Q(\buffer[8][2][4] [3]), .QN());
   DFF_X1 \buffer_reg[8][2][4][2]  (.D(\input_filter[2][4] [2]), .CK(n_55_4), 
      .Q(\buffer[8][2][4] [2]), .QN());
   DFF_X1 \buffer_reg[8][2][4][1]  (.D(\input_filter[2][4] [1]), .CK(n_55_4), 
      .Q(\buffer[8][2][4] [1]), .QN());
   DFF_X1 \buffer_reg[8][2][4][0]  (.D(\input_filter[2][4] [0]), .CK(n_55_4), 
      .Q(\buffer[8][2][4] [0]), .QN());
   DFF_X1 \buffer_reg[7][2][4][15]  (.D(\input_filter[2][4] [15]), .CK(n_55_5), 
      .Q(\buffer[7][2][4] [15]), .QN());
   DFF_X1 \buffer_reg[7][2][4][14]  (.D(\input_filter[2][4] [14]), .CK(n_55_5), 
      .Q(\buffer[7][2][4] [14]), .QN());
   DFF_X1 \buffer_reg[7][2][4][13]  (.D(\input_filter[2][4] [13]), .CK(n_55_5), 
      .Q(\buffer[7][2][4] [13]), .QN());
   DFF_X1 \buffer_reg[7][2][4][12]  (.D(\input_filter[2][4] [12]), .CK(n_55_5), 
      .Q(\buffer[7][2][4] [12]), .QN());
   DFF_X1 \buffer_reg[7][2][4][11]  (.D(\input_filter[2][4] [11]), .CK(n_55_5), 
      .Q(\buffer[7][2][4] [11]), .QN());
   DFF_X1 \buffer_reg[7][2][4][10]  (.D(\input_filter[2][4] [10]), .CK(n_55_5), 
      .Q(\buffer[7][2][4] [10]), .QN());
   DFF_X1 \buffer_reg[7][2][4][9]  (.D(\input_filter[2][4] [9]), .CK(n_55_5), 
      .Q(\buffer[7][2][4] [9]), .QN());
   DFF_X1 \buffer_reg[7][2][4][8]  (.D(\input_filter[2][4] [8]), .CK(n_55_5), 
      .Q(\buffer[7][2][4] [8]), .QN());
   DFF_X1 \buffer_reg[7][2][4][7]  (.D(\input_filter[2][4] [7]), .CK(n_55_5), 
      .Q(\buffer[7][2][4] [7]), .QN());
   DFF_X1 \buffer_reg[7][2][4][6]  (.D(\input_filter[2][4] [6]), .CK(n_55_5), 
      .Q(\buffer[7][2][4] [6]), .QN());
   DFF_X1 \buffer_reg[7][2][4][5]  (.D(\input_filter[2][4] [5]), .CK(n_55_5), 
      .Q(\buffer[7][2][4] [5]), .QN());
   DFF_X1 \buffer_reg[7][2][4][4]  (.D(\input_filter[2][4] [4]), .CK(n_55_5), 
      .Q(\buffer[7][2][4] [4]), .QN());
   DFF_X1 \buffer_reg[7][2][4][3]  (.D(\input_filter[2][4] [3]), .CK(n_55_5), 
      .Q(\buffer[7][2][4] [3]), .QN());
   DFF_X1 \buffer_reg[7][2][4][2]  (.D(\input_filter[2][4] [2]), .CK(n_55_5), 
      .Q(\buffer[7][2][4] [2]), .QN());
   DFF_X1 \buffer_reg[7][2][4][1]  (.D(\input_filter[2][4] [1]), .CK(n_55_5), 
      .Q(\buffer[7][2][4] [1]), .QN());
   DFF_X1 \buffer_reg[7][2][4][0]  (.D(\input_filter[2][4] [0]), .CK(n_55_5), 
      .Q(\buffer[7][2][4] [0]), .QN());
   DFF_X1 \buffer_reg[6][2][4][15]  (.D(\input_filter[2][4] [15]), .CK(n_55_6), 
      .Q(\buffer[6][2][4] [15]), .QN());
   DFF_X1 \buffer_reg[6][2][4][14]  (.D(\input_filter[2][4] [14]), .CK(n_55_6), 
      .Q(\buffer[6][2][4] [14]), .QN());
   DFF_X1 \buffer_reg[6][2][4][13]  (.D(\input_filter[2][4] [13]), .CK(n_55_6), 
      .Q(\buffer[6][2][4] [13]), .QN());
   DFF_X1 \buffer_reg[6][2][4][12]  (.D(\input_filter[2][4] [12]), .CK(n_55_6), 
      .Q(\buffer[6][2][4] [12]), .QN());
   DFF_X1 \buffer_reg[6][2][4][11]  (.D(\input_filter[2][4] [11]), .CK(n_55_6), 
      .Q(\buffer[6][2][4] [11]), .QN());
   DFF_X1 \buffer_reg[6][2][4][10]  (.D(\input_filter[2][4] [10]), .CK(n_55_6), 
      .Q(\buffer[6][2][4] [10]), .QN());
   DFF_X1 \buffer_reg[6][2][4][9]  (.D(\input_filter[2][4] [9]), .CK(n_55_6), 
      .Q(\buffer[6][2][4] [9]), .QN());
   DFF_X1 \buffer_reg[6][2][4][8]  (.D(\input_filter[2][4] [8]), .CK(n_55_6), 
      .Q(\buffer[6][2][4] [8]), .QN());
   DFF_X1 \buffer_reg[6][2][4][7]  (.D(\input_filter[2][4] [7]), .CK(n_55_6), 
      .Q(\buffer[6][2][4] [7]), .QN());
   DFF_X1 \buffer_reg[6][2][4][6]  (.D(\input_filter[2][4] [6]), .CK(n_55_6), 
      .Q(\buffer[6][2][4] [6]), .QN());
   DFF_X1 \buffer_reg[6][2][4][5]  (.D(\input_filter[2][4] [5]), .CK(n_55_6), 
      .Q(\buffer[6][2][4] [5]), .QN());
   DFF_X1 \buffer_reg[6][2][4][4]  (.D(\input_filter[2][4] [4]), .CK(n_55_6), 
      .Q(\buffer[6][2][4] [4]), .QN());
   DFF_X1 \buffer_reg[6][2][4][3]  (.D(\input_filter[2][4] [3]), .CK(n_55_6), 
      .Q(\buffer[6][2][4] [3]), .QN());
   DFF_X1 \buffer_reg[6][2][4][2]  (.D(\input_filter[2][4] [2]), .CK(n_55_6), 
      .Q(\buffer[6][2][4] [2]), .QN());
   DFF_X1 \buffer_reg[6][2][4][1]  (.D(\input_filter[2][4] [1]), .CK(n_55_6), 
      .Q(\buffer[6][2][4] [1]), .QN());
   DFF_X1 \buffer_reg[6][2][4][0]  (.D(\input_filter[2][4] [0]), .CK(n_55_6), 
      .Q(\buffer[6][2][4] [0]), .QN());
   DFF_X1 \buffer_reg[5][2][4][15]  (.D(\input_filter[2][4] [15]), .CK(n_55_7), 
      .Q(\buffer[5][2][4] [15]), .QN());
   DFF_X1 \buffer_reg[5][2][4][14]  (.D(\input_filter[2][4] [14]), .CK(n_55_7), 
      .Q(\buffer[5][2][4] [14]), .QN());
   DFF_X1 \buffer_reg[5][2][4][13]  (.D(\input_filter[2][4] [13]), .CK(n_55_7), 
      .Q(\buffer[5][2][4] [13]), .QN());
   DFF_X1 \buffer_reg[5][2][4][12]  (.D(\input_filter[2][4] [12]), .CK(n_55_7), 
      .Q(\buffer[5][2][4] [12]), .QN());
   DFF_X1 \buffer_reg[5][2][4][11]  (.D(\input_filter[2][4] [11]), .CK(n_55_7), 
      .Q(\buffer[5][2][4] [11]), .QN());
   DFF_X1 \buffer_reg[5][2][4][10]  (.D(\input_filter[2][4] [10]), .CK(n_55_7), 
      .Q(\buffer[5][2][4] [10]), .QN());
   DFF_X1 \buffer_reg[5][2][4][9]  (.D(\input_filter[2][4] [9]), .CK(n_55_7), 
      .Q(\buffer[5][2][4] [9]), .QN());
   DFF_X1 \buffer_reg[5][2][4][8]  (.D(\input_filter[2][4] [8]), .CK(n_55_7), 
      .Q(\buffer[5][2][4] [8]), .QN());
   DFF_X1 \buffer_reg[5][2][4][7]  (.D(\input_filter[2][4] [7]), .CK(n_55_7), 
      .Q(\buffer[5][2][4] [7]), .QN());
   DFF_X1 \buffer_reg[5][2][4][6]  (.D(\input_filter[2][4] [6]), .CK(n_55_7), 
      .Q(\buffer[5][2][4] [6]), .QN());
   DFF_X1 \buffer_reg[5][2][4][5]  (.D(\input_filter[2][4] [5]), .CK(n_55_7), 
      .Q(\buffer[5][2][4] [5]), .QN());
   DFF_X1 \buffer_reg[5][2][4][4]  (.D(\input_filter[2][4] [4]), .CK(n_55_7), 
      .Q(\buffer[5][2][4] [4]), .QN());
   DFF_X1 \buffer_reg[5][2][4][3]  (.D(\input_filter[2][4] [3]), .CK(n_55_7), 
      .Q(\buffer[5][2][4] [3]), .QN());
   DFF_X1 \buffer_reg[5][2][4][2]  (.D(\input_filter[2][4] [2]), .CK(n_55_7), 
      .Q(\buffer[5][2][4] [2]), .QN());
   DFF_X1 \buffer_reg[5][2][4][1]  (.D(\input_filter[2][4] [1]), .CK(n_55_7), 
      .Q(\buffer[5][2][4] [1]), .QN());
   DFF_X1 \buffer_reg[5][2][4][0]  (.D(\input_filter[2][4] [0]), .CK(n_55_7), 
      .Q(\buffer[5][2][4] [0]), .QN());
   DFF_X1 \buffer_reg[4][2][4][15]  (.D(\input_filter[2][4] [15]), .CK(n_55_8), 
      .Q(\buffer[4][2][4] [15]), .QN());
   DFF_X1 \buffer_reg[4][2][4][14]  (.D(\input_filter[2][4] [14]), .CK(n_55_8), 
      .Q(\buffer[4][2][4] [14]), .QN());
   DFF_X1 \buffer_reg[4][2][4][13]  (.D(\input_filter[2][4] [13]), .CK(n_55_8), 
      .Q(\buffer[4][2][4] [13]), .QN());
   DFF_X1 \buffer_reg[4][2][4][12]  (.D(\input_filter[2][4] [12]), .CK(n_55_8), 
      .Q(\buffer[4][2][4] [12]), .QN());
   DFF_X1 \buffer_reg[4][2][4][11]  (.D(\input_filter[2][4] [11]), .CK(n_55_8), 
      .Q(\buffer[4][2][4] [11]), .QN());
   DFF_X1 \buffer_reg[4][2][4][10]  (.D(\input_filter[2][4] [10]), .CK(n_55_8), 
      .Q(\buffer[4][2][4] [10]), .QN());
   DFF_X1 \buffer_reg[4][2][4][9]  (.D(\input_filter[2][4] [9]), .CK(n_55_8), 
      .Q(\buffer[4][2][4] [9]), .QN());
   DFF_X1 \buffer_reg[4][2][4][8]  (.D(\input_filter[2][4] [8]), .CK(n_55_8), 
      .Q(\buffer[4][2][4] [8]), .QN());
   DFF_X1 \buffer_reg[4][2][4][7]  (.D(\input_filter[2][4] [7]), .CK(n_55_8), 
      .Q(\buffer[4][2][4] [7]), .QN());
   DFF_X1 \buffer_reg[4][2][4][6]  (.D(\input_filter[2][4] [6]), .CK(n_55_8), 
      .Q(\buffer[4][2][4] [6]), .QN());
   DFF_X1 \buffer_reg[4][2][4][5]  (.D(\input_filter[2][4] [5]), .CK(n_55_8), 
      .Q(\buffer[4][2][4] [5]), .QN());
   DFF_X1 \buffer_reg[4][2][4][4]  (.D(\input_filter[2][4] [4]), .CK(n_55_8), 
      .Q(\buffer[4][2][4] [4]), .QN());
   DFF_X1 \buffer_reg[4][2][4][3]  (.D(\input_filter[2][4] [3]), .CK(n_55_8), 
      .Q(\buffer[4][2][4] [3]), .QN());
   DFF_X1 \buffer_reg[4][2][4][2]  (.D(\input_filter[2][4] [2]), .CK(n_55_8), 
      .Q(\buffer[4][2][4] [2]), .QN());
   DFF_X1 \buffer_reg[4][2][4][1]  (.D(\input_filter[2][4] [1]), .CK(n_55_8), 
      .Q(\buffer[4][2][4] [1]), .QN());
   DFF_X1 \buffer_reg[4][2][4][0]  (.D(\input_filter[2][4] [0]), .CK(n_55_8), 
      .Q(\buffer[4][2][4] [0]), .QN());
   DFF_X1 \buffer_reg[3][2][4][15]  (.D(\input_filter[2][4] [15]), .CK(n_55_9), 
      .Q(\buffer[3][2][4] [15]), .QN());
   DFF_X1 \buffer_reg[3][2][4][14]  (.D(\input_filter[2][4] [14]), .CK(n_55_9), 
      .Q(\buffer[3][2][4] [14]), .QN());
   DFF_X1 \buffer_reg[3][2][4][13]  (.D(\input_filter[2][4] [13]), .CK(n_55_9), 
      .Q(\buffer[3][2][4] [13]), .QN());
   DFF_X1 \buffer_reg[3][2][4][12]  (.D(\input_filter[2][4] [12]), .CK(n_55_9), 
      .Q(\buffer[3][2][4] [12]), .QN());
   DFF_X1 \buffer_reg[3][2][4][11]  (.D(\input_filter[2][4] [11]), .CK(n_55_9), 
      .Q(\buffer[3][2][4] [11]), .QN());
   DFF_X1 \buffer_reg[3][2][4][10]  (.D(\input_filter[2][4] [10]), .CK(n_55_9), 
      .Q(\buffer[3][2][4] [10]), .QN());
   DFF_X1 \buffer_reg[3][2][4][9]  (.D(\input_filter[2][4] [9]), .CK(n_55_9), 
      .Q(\buffer[3][2][4] [9]), .QN());
   DFF_X1 \buffer_reg[3][2][4][8]  (.D(\input_filter[2][4] [8]), .CK(n_55_9), 
      .Q(\buffer[3][2][4] [8]), .QN());
   DFF_X1 \buffer_reg[3][2][4][7]  (.D(\input_filter[2][4] [7]), .CK(n_55_9), 
      .Q(\buffer[3][2][4] [7]), .QN());
   DFF_X1 \buffer_reg[3][2][4][6]  (.D(\input_filter[2][4] [6]), .CK(n_55_9), 
      .Q(\buffer[3][2][4] [6]), .QN());
   DFF_X1 \buffer_reg[3][2][4][5]  (.D(\input_filter[2][4] [5]), .CK(n_55_9), 
      .Q(\buffer[3][2][4] [5]), .QN());
   DFF_X1 \buffer_reg[3][2][4][4]  (.D(\input_filter[2][4] [4]), .CK(n_55_9), 
      .Q(\buffer[3][2][4] [4]), .QN());
   DFF_X1 \buffer_reg[3][2][4][3]  (.D(\input_filter[2][4] [3]), .CK(n_55_9), 
      .Q(\buffer[3][2][4] [3]), .QN());
   DFF_X1 \buffer_reg[3][2][4][2]  (.D(\input_filter[2][4] [2]), .CK(n_55_9), 
      .Q(\buffer[3][2][4] [2]), .QN());
   DFF_X1 \buffer_reg[3][2][4][1]  (.D(\input_filter[2][4] [1]), .CK(n_55_9), 
      .Q(\buffer[3][2][4] [1]), .QN());
   DFF_X1 \buffer_reg[3][2][4][0]  (.D(\input_filter[2][4] [0]), .CK(n_55_9), 
      .Q(\buffer[3][2][4] [0]), .QN());
   DFF_X1 \buffer_reg[2][2][4][15]  (.D(\input_filter[2][4] [15]), .CK(n_55_10), 
      .Q(\buffer[2][2][4] [15]), .QN());
   DFF_X1 \buffer_reg[2][2][4][14]  (.D(\input_filter[2][4] [14]), .CK(n_55_10), 
      .Q(\buffer[2][2][4] [14]), .QN());
   DFF_X1 \buffer_reg[2][2][4][13]  (.D(\input_filter[2][4] [13]), .CK(n_55_10), 
      .Q(\buffer[2][2][4] [13]), .QN());
   DFF_X1 \buffer_reg[2][2][4][12]  (.D(\input_filter[2][4] [12]), .CK(n_55_10), 
      .Q(\buffer[2][2][4] [12]), .QN());
   DFF_X1 \buffer_reg[2][2][4][11]  (.D(\input_filter[2][4] [11]), .CK(n_55_10), 
      .Q(\buffer[2][2][4] [11]), .QN());
   DFF_X1 \buffer_reg[2][2][4][10]  (.D(\input_filter[2][4] [10]), .CK(n_55_10), 
      .Q(\buffer[2][2][4] [10]), .QN());
   DFF_X1 \buffer_reg[2][2][4][9]  (.D(\input_filter[2][4] [9]), .CK(n_55_10), 
      .Q(\buffer[2][2][4] [9]), .QN());
   DFF_X1 \buffer_reg[2][2][4][8]  (.D(\input_filter[2][4] [8]), .CK(n_55_10), 
      .Q(\buffer[2][2][4] [8]), .QN());
   DFF_X1 \buffer_reg[2][2][4][7]  (.D(\input_filter[2][4] [7]), .CK(n_55_10), 
      .Q(\buffer[2][2][4] [7]), .QN());
   DFF_X1 \buffer_reg[2][2][4][6]  (.D(\input_filter[2][4] [6]), .CK(n_55_10), 
      .Q(\buffer[2][2][4] [6]), .QN());
   DFF_X1 \buffer_reg[2][2][4][5]  (.D(\input_filter[2][4] [5]), .CK(n_55_10), 
      .Q(\buffer[2][2][4] [5]), .QN());
   DFF_X1 \buffer_reg[2][2][4][4]  (.D(\input_filter[2][4] [4]), .CK(n_55_10), 
      .Q(\buffer[2][2][4] [4]), .QN());
   DFF_X1 \buffer_reg[2][2][4][3]  (.D(\input_filter[2][4] [3]), .CK(n_55_10), 
      .Q(\buffer[2][2][4] [3]), .QN());
   DFF_X1 \buffer_reg[2][2][4][2]  (.D(\input_filter[2][4] [2]), .CK(n_55_10), 
      .Q(\buffer[2][2][4] [2]), .QN());
   DFF_X1 \buffer_reg[2][2][4][1]  (.D(\input_filter[2][4] [1]), .CK(n_55_10), 
      .Q(\buffer[2][2][4] [1]), .QN());
   DFF_X1 \buffer_reg[2][2][4][0]  (.D(\input_filter[2][4] [0]), .CK(n_55_10), 
      .Q(\buffer[2][2][4] [0]), .QN());
   DFF_X1 \buffer_reg[1][2][4][15]  (.D(\input_filter[2][4] [15]), .CK(n_55_11), 
      .Q(\buffer[1][2][4] [15]), .QN());
   DFF_X1 \buffer_reg[1][2][4][14]  (.D(\input_filter[2][4] [14]), .CK(n_55_11), 
      .Q(\buffer[1][2][4] [14]), .QN());
   DFF_X1 \buffer_reg[1][2][4][13]  (.D(\input_filter[2][4] [13]), .CK(n_55_11), 
      .Q(\buffer[1][2][4] [13]), .QN());
   DFF_X1 \buffer_reg[1][2][4][12]  (.D(\input_filter[2][4] [12]), .CK(n_55_11), 
      .Q(\buffer[1][2][4] [12]), .QN());
   DFF_X1 \buffer_reg[1][2][4][11]  (.D(\input_filter[2][4] [11]), .CK(n_55_11), 
      .Q(\buffer[1][2][4] [11]), .QN());
   DFF_X1 \buffer_reg[1][2][4][10]  (.D(\input_filter[2][4] [10]), .CK(n_55_11), 
      .Q(\buffer[1][2][4] [10]), .QN());
   DFF_X1 \buffer_reg[1][2][4][9]  (.D(\input_filter[2][4] [9]), .CK(n_55_11), 
      .Q(\buffer[1][2][4] [9]), .QN());
   DFF_X1 \buffer_reg[1][2][4][8]  (.D(\input_filter[2][4] [8]), .CK(n_55_11), 
      .Q(\buffer[1][2][4] [8]), .QN());
   DFF_X1 \buffer_reg[1][2][4][7]  (.D(\input_filter[2][4] [7]), .CK(n_55_11), 
      .Q(\buffer[1][2][4] [7]), .QN());
   DFF_X1 \buffer_reg[1][2][4][6]  (.D(\input_filter[2][4] [6]), .CK(n_55_11), 
      .Q(\buffer[1][2][4] [6]), .QN());
   DFF_X1 \buffer_reg[1][2][4][5]  (.D(\input_filter[2][4] [5]), .CK(n_55_11), 
      .Q(\buffer[1][2][4] [5]), .QN());
   DFF_X1 \buffer_reg[1][2][4][4]  (.D(\input_filter[2][4] [4]), .CK(n_55_11), 
      .Q(\buffer[1][2][4] [4]), .QN());
   DFF_X1 \buffer_reg[1][2][4][3]  (.D(\input_filter[2][4] [3]), .CK(n_55_11), 
      .Q(\buffer[1][2][4] [3]), .QN());
   DFF_X1 \buffer_reg[1][2][4][2]  (.D(\input_filter[2][4] [2]), .CK(n_55_11), 
      .Q(\buffer[1][2][4] [2]), .QN());
   DFF_X1 \buffer_reg[1][2][4][1]  (.D(\input_filter[2][4] [1]), .CK(n_55_11), 
      .Q(\buffer[1][2][4] [1]), .QN());
   DFF_X1 \buffer_reg[1][2][4][0]  (.D(\input_filter[2][4] [0]), .CK(n_55_11), 
      .Q(\buffer[1][2][4] [0]), .QN());
   DFF_X1 \buffer_reg[0][2][4][15]  (.D(\input_filter[2][4] [15]), .CK(n_55_12), 
      .Q(\buffer[0][2][4] [15]), .QN());
   DFF_X1 \buffer_reg[0][2][4][14]  (.D(\input_filter[2][4] [14]), .CK(n_55_12), 
      .Q(\buffer[0][2][4] [14]), .QN());
   DFF_X1 \buffer_reg[0][2][4][13]  (.D(\input_filter[2][4] [13]), .CK(n_55_12), 
      .Q(\buffer[0][2][4] [13]), .QN());
   DFF_X1 \buffer_reg[0][2][4][12]  (.D(\input_filter[2][4] [12]), .CK(n_55_12), 
      .Q(\buffer[0][2][4] [12]), .QN());
   DFF_X1 \buffer_reg[0][2][4][11]  (.D(\input_filter[2][4] [11]), .CK(n_55_12), 
      .Q(\buffer[0][2][4] [11]), .QN());
   DFF_X1 \buffer_reg[0][2][4][10]  (.D(\input_filter[2][4] [10]), .CK(n_55_12), 
      .Q(\buffer[0][2][4] [10]), .QN());
   DFF_X1 \buffer_reg[0][2][4][9]  (.D(\input_filter[2][4] [9]), .CK(n_55_12), 
      .Q(\buffer[0][2][4] [9]), .QN());
   DFF_X1 \buffer_reg[0][2][4][8]  (.D(\input_filter[2][4] [8]), .CK(n_55_12), 
      .Q(\buffer[0][2][4] [8]), .QN());
   DFF_X1 \buffer_reg[0][2][4][7]  (.D(\input_filter[2][4] [7]), .CK(n_55_12), 
      .Q(\buffer[0][2][4] [7]), .QN());
   DFF_X1 \buffer_reg[0][2][4][6]  (.D(\input_filter[2][4] [6]), .CK(n_55_12), 
      .Q(\buffer[0][2][4] [6]), .QN());
   DFF_X1 \buffer_reg[0][2][4][5]  (.D(\input_filter[2][4] [5]), .CK(n_55_12), 
      .Q(\buffer[0][2][4] [5]), .QN());
   DFF_X1 \buffer_reg[0][2][4][4]  (.D(\input_filter[2][4] [4]), .CK(n_55_12), 
      .Q(\buffer[0][2][4] [4]), .QN());
   DFF_X1 \buffer_reg[0][2][4][3]  (.D(\input_filter[2][4] [3]), .CK(n_55_12), 
      .Q(\buffer[0][2][4] [3]), .QN());
   DFF_X1 \buffer_reg[0][2][4][2]  (.D(\input_filter[2][4] [2]), .CK(n_55_12), 
      .Q(\buffer[0][2][4] [2]), .QN());
   DFF_X1 \buffer_reg[0][2][4][1]  (.D(\input_filter[2][4] [1]), .CK(n_55_12), 
      .Q(\buffer[0][2][4] [1]), .QN());
   DFF_X1 \buffer_reg[0][2][4][0]  (.D(\input_filter[2][4] [0]), .CK(n_55_12), 
      .Q(\buffer[0][2][4] [0]), .QN());
   DFF_X1 \buffer_reg[15][2][3][15]  (.D(\input_filter[2][3] [15]), .CK(n_55_13), 
      .Q(\buffer[15][2][3] [15]), .QN());
   DFF_X1 \buffer_reg[15][2][3][14]  (.D(\input_filter[2][3] [14]), .CK(n_55_13), 
      .Q(\buffer[15][2][3] [14]), .QN());
   DFF_X1 \buffer_reg[15][2][3][13]  (.D(\input_filter[2][3] [13]), .CK(n_55_13), 
      .Q(\buffer[15][2][3] [13]), .QN());
   DFF_X1 \buffer_reg[15][2][3][12]  (.D(\input_filter[2][3] [12]), .CK(n_55_13), 
      .Q(\buffer[15][2][3] [12]), .QN());
   DFF_X1 \buffer_reg[15][2][3][11]  (.D(\input_filter[2][3] [11]), .CK(n_55_13), 
      .Q(\buffer[15][2][3] [11]), .QN());
   DFF_X1 \buffer_reg[15][2][3][10]  (.D(\input_filter[2][3] [10]), .CK(n_55_13), 
      .Q(\buffer[15][2][3] [10]), .QN());
   DFF_X1 \buffer_reg[15][2][3][9]  (.D(\input_filter[2][3] [9]), .CK(n_55_13), 
      .Q(\buffer[15][2][3] [9]), .QN());
   DFF_X1 \buffer_reg[15][2][3][8]  (.D(\input_filter[2][3] [8]), .CK(n_55_13), 
      .Q(\buffer[15][2][3] [8]), .QN());
   DFF_X1 \buffer_reg[15][2][3][7]  (.D(\input_filter[2][3] [7]), .CK(n_55_13), 
      .Q(\buffer[15][2][3] [7]), .QN());
   DFF_X1 \buffer_reg[15][2][3][6]  (.D(\input_filter[2][3] [6]), .CK(n_55_13), 
      .Q(\buffer[15][2][3] [6]), .QN());
   DFF_X1 \buffer_reg[15][2][3][5]  (.D(\input_filter[2][3] [5]), .CK(n_55_13), 
      .Q(\buffer[15][2][3] [5]), .QN());
   DFF_X1 \buffer_reg[15][2][3][4]  (.D(\input_filter[2][3] [4]), .CK(n_55_13), 
      .Q(\buffer[15][2][3] [4]), .QN());
   DFF_X1 \buffer_reg[15][2][3][3]  (.D(\input_filter[2][3] [3]), .CK(n_55_13), 
      .Q(\buffer[15][2][3] [3]), .QN());
   DFF_X1 \buffer_reg[15][2][3][2]  (.D(\input_filter[2][3] [2]), .CK(n_55_13), 
      .Q(\buffer[15][2][3] [2]), .QN());
   DFF_X1 \buffer_reg[15][2][3][1]  (.D(\input_filter[2][3] [1]), .CK(n_55_13), 
      .Q(\buffer[15][2][3] [1]), .QN());
   DFF_X1 \buffer_reg[15][2][3][0]  (.D(\input_filter[2][3] [0]), .CK(n_55_13), 
      .Q(\buffer[15][2][3] [0]), .QN());
   DFF_X1 \buffer_reg[14][2][3][15]  (.D(\input_filter[2][3] [15]), .CK(n_55_14), 
      .Q(\buffer[14][2][3] [15]), .QN());
   DFF_X1 \buffer_reg[14][2][3][14]  (.D(\input_filter[2][3] [14]), .CK(n_55_14), 
      .Q(\buffer[14][2][3] [14]), .QN());
   DFF_X1 \buffer_reg[14][2][3][13]  (.D(\input_filter[2][3] [13]), .CK(n_55_14), 
      .Q(\buffer[14][2][3] [13]), .QN());
   DFF_X1 \buffer_reg[14][2][3][12]  (.D(\input_filter[2][3] [12]), .CK(n_55_14), 
      .Q(\buffer[14][2][3] [12]), .QN());
   DFF_X1 \buffer_reg[14][2][3][11]  (.D(\input_filter[2][3] [11]), .CK(n_55_14), 
      .Q(\buffer[14][2][3] [11]), .QN());
   DFF_X1 \buffer_reg[14][2][3][10]  (.D(\input_filter[2][3] [10]), .CK(n_55_14), 
      .Q(\buffer[14][2][3] [10]), .QN());
   DFF_X1 \buffer_reg[14][2][3][9]  (.D(\input_filter[2][3] [9]), .CK(n_55_14), 
      .Q(\buffer[14][2][3] [9]), .QN());
   DFF_X1 \buffer_reg[14][2][3][8]  (.D(\input_filter[2][3] [8]), .CK(n_55_14), 
      .Q(\buffer[14][2][3] [8]), .QN());
   DFF_X1 \buffer_reg[14][2][3][7]  (.D(\input_filter[2][3] [7]), .CK(n_55_14), 
      .Q(\buffer[14][2][3] [7]), .QN());
   DFF_X1 \buffer_reg[14][2][3][6]  (.D(\input_filter[2][3] [6]), .CK(n_55_14), 
      .Q(\buffer[14][2][3] [6]), .QN());
   DFF_X1 \buffer_reg[14][2][3][5]  (.D(\input_filter[2][3] [5]), .CK(n_55_14), 
      .Q(\buffer[14][2][3] [5]), .QN());
   DFF_X1 \buffer_reg[14][2][3][4]  (.D(\input_filter[2][3] [4]), .CK(n_55_14), 
      .Q(\buffer[14][2][3] [4]), .QN());
   DFF_X1 \buffer_reg[14][2][3][3]  (.D(\input_filter[2][3] [3]), .CK(n_55_14), 
      .Q(\buffer[14][2][3] [3]), .QN());
   DFF_X1 \buffer_reg[14][2][3][2]  (.D(\input_filter[2][3] [2]), .CK(n_55_14), 
      .Q(\buffer[14][2][3] [2]), .QN());
   DFF_X1 \buffer_reg[14][2][3][1]  (.D(\input_filter[2][3] [1]), .CK(n_55_14), 
      .Q(\buffer[14][2][3] [1]), .QN());
   DFF_X1 \buffer_reg[14][2][3][0]  (.D(\input_filter[2][3] [0]), .CK(n_55_14), 
      .Q(\buffer[14][2][3] [0]), .QN());
   DFF_X1 \buffer_reg[13][2][3][15]  (.D(\input_filter[2][3] [15]), .CK(n_55_15), 
      .Q(\buffer[13][2][3] [15]), .QN());
   DFF_X1 \buffer_reg[13][2][3][14]  (.D(\input_filter[2][3] [14]), .CK(n_55_15), 
      .Q(\buffer[13][2][3] [14]), .QN());
   DFF_X1 \buffer_reg[13][2][3][13]  (.D(\input_filter[2][3] [13]), .CK(n_55_15), 
      .Q(\buffer[13][2][3] [13]), .QN());
   DFF_X1 \buffer_reg[13][2][3][12]  (.D(\input_filter[2][3] [12]), .CK(n_55_15), 
      .Q(\buffer[13][2][3] [12]), .QN());
   DFF_X1 \buffer_reg[13][2][3][11]  (.D(\input_filter[2][3] [11]), .CK(n_55_15), 
      .Q(\buffer[13][2][3] [11]), .QN());
   DFF_X1 \buffer_reg[13][2][3][10]  (.D(\input_filter[2][3] [10]), .CK(n_55_15), 
      .Q(\buffer[13][2][3] [10]), .QN());
   DFF_X1 \buffer_reg[13][2][3][9]  (.D(\input_filter[2][3] [9]), .CK(n_55_15), 
      .Q(\buffer[13][2][3] [9]), .QN());
   DFF_X1 \buffer_reg[13][2][3][8]  (.D(\input_filter[2][3] [8]), .CK(n_55_15), 
      .Q(\buffer[13][2][3] [8]), .QN());
   DFF_X1 \buffer_reg[13][2][3][7]  (.D(\input_filter[2][3] [7]), .CK(n_55_15), 
      .Q(\buffer[13][2][3] [7]), .QN());
   DFF_X1 \buffer_reg[13][2][3][6]  (.D(\input_filter[2][3] [6]), .CK(n_55_15), 
      .Q(\buffer[13][2][3] [6]), .QN());
   DFF_X1 \buffer_reg[13][2][3][5]  (.D(\input_filter[2][3] [5]), .CK(n_55_15), 
      .Q(\buffer[13][2][3] [5]), .QN());
   DFF_X1 \buffer_reg[13][2][3][4]  (.D(\input_filter[2][3] [4]), .CK(n_55_15), 
      .Q(\buffer[13][2][3] [4]), .QN());
   DFF_X1 \buffer_reg[13][2][3][3]  (.D(\input_filter[2][3] [3]), .CK(n_55_15), 
      .Q(\buffer[13][2][3] [3]), .QN());
   DFF_X1 \buffer_reg[13][2][3][2]  (.D(\input_filter[2][3] [2]), .CK(n_55_15), 
      .Q(\buffer[13][2][3] [2]), .QN());
   DFF_X1 \buffer_reg[13][2][3][1]  (.D(\input_filter[2][3] [1]), .CK(n_55_15), 
      .Q(\buffer[13][2][3] [1]), .QN());
   DFF_X1 \buffer_reg[13][2][3][0]  (.D(\input_filter[2][3] [0]), .CK(n_55_15), 
      .Q(\buffer[13][2][3] [0]), .QN());
   DFF_X1 \buffer_reg[12][2][3][15]  (.D(\input_filter[2][3] [15]), .CK(n_55_0), 
      .Q(\buffer[12][2][3] [15]), .QN());
   DFF_X1 \buffer_reg[12][2][3][14]  (.D(\input_filter[2][3] [14]), .CK(n_55_0), 
      .Q(\buffer[12][2][3] [14]), .QN());
   DFF_X1 \buffer_reg[12][2][3][13]  (.D(\input_filter[2][3] [13]), .CK(n_55_0), 
      .Q(\buffer[12][2][3] [13]), .QN());
   DFF_X1 \buffer_reg[12][2][3][12]  (.D(\input_filter[2][3] [12]), .CK(n_55_0), 
      .Q(\buffer[12][2][3] [12]), .QN());
   DFF_X1 \buffer_reg[12][2][3][11]  (.D(\input_filter[2][3] [11]), .CK(n_55_0), 
      .Q(\buffer[12][2][3] [11]), .QN());
   DFF_X1 \buffer_reg[12][2][3][10]  (.D(\input_filter[2][3] [10]), .CK(n_55_0), 
      .Q(\buffer[12][2][3] [10]), .QN());
   DFF_X1 \buffer_reg[12][2][3][9]  (.D(\input_filter[2][3] [9]), .CK(n_55_0), 
      .Q(\buffer[12][2][3] [9]), .QN());
   DFF_X1 \buffer_reg[12][2][3][8]  (.D(\input_filter[2][3] [8]), .CK(n_55_0), 
      .Q(\buffer[12][2][3] [8]), .QN());
   DFF_X1 \buffer_reg[12][2][3][7]  (.D(\input_filter[2][3] [7]), .CK(n_55_0), 
      .Q(\buffer[12][2][3] [7]), .QN());
   DFF_X1 \buffer_reg[12][2][3][6]  (.D(\input_filter[2][3] [6]), .CK(n_55_0), 
      .Q(\buffer[12][2][3] [6]), .QN());
   DFF_X1 \buffer_reg[12][2][3][5]  (.D(\input_filter[2][3] [5]), .CK(n_55_0), 
      .Q(\buffer[12][2][3] [5]), .QN());
   DFF_X1 \buffer_reg[12][2][3][4]  (.D(\input_filter[2][3] [4]), .CK(n_55_0), 
      .Q(\buffer[12][2][3] [4]), .QN());
   DFF_X1 \buffer_reg[12][2][3][3]  (.D(\input_filter[2][3] [3]), .CK(n_55_0), 
      .Q(\buffer[12][2][3] [3]), .QN());
   DFF_X1 \buffer_reg[12][2][3][2]  (.D(\input_filter[2][3] [2]), .CK(n_55_0), 
      .Q(\buffer[12][2][3] [2]), .QN());
   DFF_X1 \buffer_reg[12][2][3][1]  (.D(\input_filter[2][3] [1]), .CK(n_55_0), 
      .Q(\buffer[12][2][3] [1]), .QN());
   DFF_X1 \buffer_reg[12][2][3][0]  (.D(\input_filter[2][3] [0]), .CK(n_55_0), 
      .Q(\buffer[12][2][3] [0]), .QN());
   DFF_X1 \buffer_reg[11][2][3][15]  (.D(\input_filter[2][3] [15]), .CK(n_55_1), 
      .Q(\buffer[11][2][3] [15]), .QN());
   DFF_X1 \buffer_reg[11][2][3][14]  (.D(\input_filter[2][3] [14]), .CK(n_55_1), 
      .Q(\buffer[11][2][3] [14]), .QN());
   DFF_X1 \buffer_reg[11][2][3][13]  (.D(\input_filter[2][3] [13]), .CK(n_55_1), 
      .Q(\buffer[11][2][3] [13]), .QN());
   DFF_X1 \buffer_reg[11][2][3][12]  (.D(\input_filter[2][3] [12]), .CK(n_55_1), 
      .Q(\buffer[11][2][3] [12]), .QN());
   DFF_X1 \buffer_reg[11][2][3][11]  (.D(\input_filter[2][3] [11]), .CK(n_55_1), 
      .Q(\buffer[11][2][3] [11]), .QN());
   DFF_X1 \buffer_reg[11][2][3][10]  (.D(\input_filter[2][3] [10]), .CK(n_55_1), 
      .Q(\buffer[11][2][3] [10]), .QN());
   DFF_X1 \buffer_reg[11][2][3][9]  (.D(\input_filter[2][3] [9]), .CK(n_55_1), 
      .Q(\buffer[11][2][3] [9]), .QN());
   DFF_X1 \buffer_reg[11][2][3][8]  (.D(\input_filter[2][3] [8]), .CK(n_55_1), 
      .Q(\buffer[11][2][3] [8]), .QN());
   DFF_X1 \buffer_reg[11][2][3][7]  (.D(\input_filter[2][3] [7]), .CK(n_55_1), 
      .Q(\buffer[11][2][3] [7]), .QN());
   DFF_X1 \buffer_reg[11][2][3][6]  (.D(\input_filter[2][3] [6]), .CK(n_55_1), 
      .Q(\buffer[11][2][3] [6]), .QN());
   DFF_X1 \buffer_reg[11][2][3][5]  (.D(\input_filter[2][3] [5]), .CK(n_55_1), 
      .Q(\buffer[11][2][3] [5]), .QN());
   DFF_X1 \buffer_reg[11][2][3][4]  (.D(\input_filter[2][3] [4]), .CK(n_55_1), 
      .Q(\buffer[11][2][3] [4]), .QN());
   DFF_X1 \buffer_reg[11][2][3][3]  (.D(\input_filter[2][3] [3]), .CK(n_55_1), 
      .Q(\buffer[11][2][3] [3]), .QN());
   DFF_X1 \buffer_reg[11][2][3][2]  (.D(\input_filter[2][3] [2]), .CK(n_55_1), 
      .Q(\buffer[11][2][3] [2]), .QN());
   DFF_X1 \buffer_reg[11][2][3][1]  (.D(\input_filter[2][3] [1]), .CK(n_55_1), 
      .Q(\buffer[11][2][3] [1]), .QN());
   DFF_X1 \buffer_reg[11][2][3][0]  (.D(\input_filter[2][3] [0]), .CK(n_55_1), 
      .Q(\buffer[11][2][3] [0]), .QN());
   DFF_X1 \buffer_reg[10][2][3][15]  (.D(\input_filter[2][3] [15]), .CK(n_55_2), 
      .Q(\buffer[10][2][3] [15]), .QN());
   DFF_X1 \buffer_reg[10][2][3][14]  (.D(\input_filter[2][3] [14]), .CK(n_55_2), 
      .Q(\buffer[10][2][3] [14]), .QN());
   DFF_X1 \buffer_reg[10][2][3][13]  (.D(\input_filter[2][3] [13]), .CK(n_55_2), 
      .Q(\buffer[10][2][3] [13]), .QN());
   DFF_X1 \buffer_reg[10][2][3][12]  (.D(\input_filter[2][3] [12]), .CK(n_55_2), 
      .Q(\buffer[10][2][3] [12]), .QN());
   DFF_X1 \buffer_reg[10][2][3][11]  (.D(\input_filter[2][3] [11]), .CK(n_55_2), 
      .Q(\buffer[10][2][3] [11]), .QN());
   DFF_X1 \buffer_reg[10][2][3][10]  (.D(\input_filter[2][3] [10]), .CK(n_55_2), 
      .Q(\buffer[10][2][3] [10]), .QN());
   DFF_X1 \buffer_reg[10][2][3][9]  (.D(\input_filter[2][3] [9]), .CK(n_55_2), 
      .Q(\buffer[10][2][3] [9]), .QN());
   DFF_X1 \buffer_reg[10][2][3][8]  (.D(\input_filter[2][3] [8]), .CK(n_55_2), 
      .Q(\buffer[10][2][3] [8]), .QN());
   DFF_X1 \buffer_reg[10][2][3][7]  (.D(\input_filter[2][3] [7]), .CK(n_55_2), 
      .Q(\buffer[10][2][3] [7]), .QN());
   DFF_X1 \buffer_reg[10][2][3][6]  (.D(\input_filter[2][3] [6]), .CK(n_55_2), 
      .Q(\buffer[10][2][3] [6]), .QN());
   DFF_X1 \buffer_reg[10][2][3][5]  (.D(\input_filter[2][3] [5]), .CK(n_55_2), 
      .Q(\buffer[10][2][3] [5]), .QN());
   DFF_X1 \buffer_reg[10][2][3][4]  (.D(\input_filter[2][3] [4]), .CK(n_55_2), 
      .Q(\buffer[10][2][3] [4]), .QN());
   DFF_X1 \buffer_reg[10][2][3][3]  (.D(\input_filter[2][3] [3]), .CK(n_55_2), 
      .Q(\buffer[10][2][3] [3]), .QN());
   DFF_X1 \buffer_reg[10][2][3][2]  (.D(\input_filter[2][3] [2]), .CK(n_55_2), 
      .Q(\buffer[10][2][3] [2]), .QN());
   DFF_X1 \buffer_reg[10][2][3][1]  (.D(\input_filter[2][3] [1]), .CK(n_55_2), 
      .Q(\buffer[10][2][3] [1]), .QN());
   DFF_X1 \buffer_reg[10][2][3][0]  (.D(\input_filter[2][3] [0]), .CK(n_55_2), 
      .Q(\buffer[10][2][3] [0]), .QN());
   DFF_X1 \buffer_reg[9][2][3][15]  (.D(\input_filter[2][3] [15]), .CK(n_55_3), 
      .Q(\buffer[9][2][3] [15]), .QN());
   DFF_X1 \buffer_reg[9][2][3][14]  (.D(\input_filter[2][3] [14]), .CK(n_55_3), 
      .Q(\buffer[9][2][3] [14]), .QN());
   DFF_X1 \buffer_reg[9][2][3][13]  (.D(\input_filter[2][3] [13]), .CK(n_55_3), 
      .Q(\buffer[9][2][3] [13]), .QN());
   DFF_X1 \buffer_reg[9][2][3][12]  (.D(\input_filter[2][3] [12]), .CK(n_55_3), 
      .Q(\buffer[9][2][3] [12]), .QN());
   DFF_X1 \buffer_reg[9][2][3][11]  (.D(\input_filter[2][3] [11]), .CK(n_55_3), 
      .Q(\buffer[9][2][3] [11]), .QN());
   DFF_X1 \buffer_reg[9][2][3][10]  (.D(\input_filter[2][3] [10]), .CK(n_55_3), 
      .Q(\buffer[9][2][3] [10]), .QN());
   DFF_X1 \buffer_reg[9][2][3][9]  (.D(\input_filter[2][3] [9]), .CK(n_55_3), 
      .Q(\buffer[9][2][3] [9]), .QN());
   DFF_X1 \buffer_reg[9][2][3][8]  (.D(\input_filter[2][3] [8]), .CK(n_55_3), 
      .Q(\buffer[9][2][3] [8]), .QN());
   DFF_X1 \buffer_reg[9][2][3][7]  (.D(\input_filter[2][3] [7]), .CK(n_55_3), 
      .Q(\buffer[9][2][3] [7]), .QN());
   DFF_X1 \buffer_reg[9][2][3][6]  (.D(\input_filter[2][3] [6]), .CK(n_55_3), 
      .Q(\buffer[9][2][3] [6]), .QN());
   DFF_X1 \buffer_reg[9][2][3][5]  (.D(\input_filter[2][3] [5]), .CK(n_55_3), 
      .Q(\buffer[9][2][3] [5]), .QN());
   DFF_X1 \buffer_reg[9][2][3][4]  (.D(\input_filter[2][3] [4]), .CK(n_55_3), 
      .Q(\buffer[9][2][3] [4]), .QN());
   DFF_X1 \buffer_reg[9][2][3][3]  (.D(\input_filter[2][3] [3]), .CK(n_55_3), 
      .Q(\buffer[9][2][3] [3]), .QN());
   DFF_X1 \buffer_reg[9][2][3][2]  (.D(\input_filter[2][3] [2]), .CK(n_55_3), 
      .Q(\buffer[9][2][3] [2]), .QN());
   DFF_X1 \buffer_reg[9][2][3][1]  (.D(\input_filter[2][3] [1]), .CK(n_55_3), 
      .Q(\buffer[9][2][3] [1]), .QN());
   DFF_X1 \buffer_reg[9][2][3][0]  (.D(\input_filter[2][3] [0]), .CK(n_55_3), 
      .Q(\buffer[9][2][3] [0]), .QN());
   DFF_X1 \buffer_reg[8][2][3][15]  (.D(\input_filter[2][3] [15]), .CK(n_55_4), 
      .Q(\buffer[8][2][3] [15]), .QN());
   DFF_X1 \buffer_reg[8][2][3][14]  (.D(\input_filter[2][3] [14]), .CK(n_55_4), 
      .Q(\buffer[8][2][3] [14]), .QN());
   DFF_X1 \buffer_reg[8][2][3][13]  (.D(\input_filter[2][3] [13]), .CK(n_55_4), 
      .Q(\buffer[8][2][3] [13]), .QN());
   DFF_X1 \buffer_reg[8][2][3][12]  (.D(\input_filter[2][3] [12]), .CK(n_55_4), 
      .Q(\buffer[8][2][3] [12]), .QN());
   DFF_X1 \buffer_reg[8][2][3][11]  (.D(\input_filter[2][3] [11]), .CK(n_55_4), 
      .Q(\buffer[8][2][3] [11]), .QN());
   DFF_X1 \buffer_reg[8][2][3][10]  (.D(\input_filter[2][3] [10]), .CK(n_55_4), 
      .Q(\buffer[8][2][3] [10]), .QN());
   DFF_X1 \buffer_reg[8][2][3][9]  (.D(\input_filter[2][3] [9]), .CK(n_55_4), 
      .Q(\buffer[8][2][3] [9]), .QN());
   DFF_X1 \buffer_reg[8][2][3][8]  (.D(\input_filter[2][3] [8]), .CK(n_55_4), 
      .Q(\buffer[8][2][3] [8]), .QN());
   DFF_X1 \buffer_reg[8][2][3][7]  (.D(\input_filter[2][3] [7]), .CK(n_55_4), 
      .Q(\buffer[8][2][3] [7]), .QN());
   DFF_X1 \buffer_reg[8][2][3][6]  (.D(\input_filter[2][3] [6]), .CK(n_55_4), 
      .Q(\buffer[8][2][3] [6]), .QN());
   DFF_X1 \buffer_reg[8][2][3][5]  (.D(\input_filter[2][3] [5]), .CK(n_55_4), 
      .Q(\buffer[8][2][3] [5]), .QN());
   DFF_X1 \buffer_reg[8][2][3][4]  (.D(\input_filter[2][3] [4]), .CK(n_55_4), 
      .Q(\buffer[8][2][3] [4]), .QN());
   DFF_X1 \buffer_reg[8][2][3][3]  (.D(\input_filter[2][3] [3]), .CK(n_55_4), 
      .Q(\buffer[8][2][3] [3]), .QN());
   DFF_X1 \buffer_reg[8][2][3][2]  (.D(\input_filter[2][3] [2]), .CK(n_55_4), 
      .Q(\buffer[8][2][3] [2]), .QN());
   DFF_X1 \buffer_reg[8][2][3][1]  (.D(\input_filter[2][3] [1]), .CK(n_55_4), 
      .Q(\buffer[8][2][3] [1]), .QN());
   DFF_X1 \buffer_reg[8][2][3][0]  (.D(\input_filter[2][3] [0]), .CK(n_55_4), 
      .Q(\buffer[8][2][3] [0]), .QN());
   DFF_X1 \buffer_reg[7][2][3][15]  (.D(\input_filter[2][3] [15]), .CK(n_55_5), 
      .Q(\buffer[7][2][3] [15]), .QN());
   DFF_X1 \buffer_reg[7][2][3][14]  (.D(\input_filter[2][3] [14]), .CK(n_55_5), 
      .Q(\buffer[7][2][3] [14]), .QN());
   DFF_X1 \buffer_reg[7][2][3][13]  (.D(\input_filter[2][3] [13]), .CK(n_55_5), 
      .Q(\buffer[7][2][3] [13]), .QN());
   DFF_X1 \buffer_reg[7][2][3][12]  (.D(\input_filter[2][3] [12]), .CK(n_55_5), 
      .Q(\buffer[7][2][3] [12]), .QN());
   DFF_X1 \buffer_reg[7][2][3][11]  (.D(\input_filter[2][3] [11]), .CK(n_55_5), 
      .Q(\buffer[7][2][3] [11]), .QN());
   DFF_X1 \buffer_reg[7][2][3][10]  (.D(\input_filter[2][3] [10]), .CK(n_55_5), 
      .Q(\buffer[7][2][3] [10]), .QN());
   DFF_X1 \buffer_reg[7][2][3][9]  (.D(\input_filter[2][3] [9]), .CK(n_55_5), 
      .Q(\buffer[7][2][3] [9]), .QN());
   DFF_X1 \buffer_reg[7][2][3][8]  (.D(\input_filter[2][3] [8]), .CK(n_55_5), 
      .Q(\buffer[7][2][3] [8]), .QN());
   DFF_X1 \buffer_reg[7][2][3][7]  (.D(\input_filter[2][3] [7]), .CK(n_55_5), 
      .Q(\buffer[7][2][3] [7]), .QN());
   DFF_X1 \buffer_reg[7][2][3][6]  (.D(\input_filter[2][3] [6]), .CK(n_55_5), 
      .Q(\buffer[7][2][3] [6]), .QN());
   DFF_X1 \buffer_reg[7][2][3][5]  (.D(\input_filter[2][3] [5]), .CK(n_55_5), 
      .Q(\buffer[7][2][3] [5]), .QN());
   DFF_X1 \buffer_reg[7][2][3][4]  (.D(\input_filter[2][3] [4]), .CK(n_55_5), 
      .Q(\buffer[7][2][3] [4]), .QN());
   DFF_X1 \buffer_reg[7][2][3][3]  (.D(\input_filter[2][3] [3]), .CK(n_55_5), 
      .Q(\buffer[7][2][3] [3]), .QN());
   DFF_X1 \buffer_reg[7][2][3][2]  (.D(\input_filter[2][3] [2]), .CK(n_55_5), 
      .Q(\buffer[7][2][3] [2]), .QN());
   DFF_X1 \buffer_reg[7][2][3][1]  (.D(\input_filter[2][3] [1]), .CK(n_55_5), 
      .Q(\buffer[7][2][3] [1]), .QN());
   DFF_X1 \buffer_reg[7][2][3][0]  (.D(\input_filter[2][3] [0]), .CK(n_55_5), 
      .Q(\buffer[7][2][3] [0]), .QN());
   DFF_X1 \buffer_reg[6][2][3][15]  (.D(\input_filter[2][3] [15]), .CK(n_55_6), 
      .Q(\buffer[6][2][3] [15]), .QN());
   DFF_X1 \buffer_reg[6][2][3][14]  (.D(\input_filter[2][3] [14]), .CK(n_55_6), 
      .Q(\buffer[6][2][3] [14]), .QN());
   DFF_X1 \buffer_reg[6][2][3][13]  (.D(\input_filter[2][3] [13]), .CK(n_55_6), 
      .Q(\buffer[6][2][3] [13]), .QN());
   DFF_X1 \buffer_reg[6][2][3][12]  (.D(\input_filter[2][3] [12]), .CK(n_55_6), 
      .Q(\buffer[6][2][3] [12]), .QN());
   DFF_X1 \buffer_reg[6][2][3][11]  (.D(\input_filter[2][3] [11]), .CK(n_55_6), 
      .Q(\buffer[6][2][3] [11]), .QN());
   DFF_X1 \buffer_reg[6][2][3][10]  (.D(\input_filter[2][3] [10]), .CK(n_55_6), 
      .Q(\buffer[6][2][3] [10]), .QN());
   DFF_X1 \buffer_reg[6][2][3][9]  (.D(\input_filter[2][3] [9]), .CK(n_55_6), 
      .Q(\buffer[6][2][3] [9]), .QN());
   DFF_X1 \buffer_reg[6][2][3][8]  (.D(\input_filter[2][3] [8]), .CK(n_55_6), 
      .Q(\buffer[6][2][3] [8]), .QN());
   DFF_X1 \buffer_reg[6][2][3][7]  (.D(\input_filter[2][3] [7]), .CK(n_55_6), 
      .Q(\buffer[6][2][3] [7]), .QN());
   DFF_X1 \buffer_reg[6][2][3][6]  (.D(\input_filter[2][3] [6]), .CK(n_55_6), 
      .Q(\buffer[6][2][3] [6]), .QN());
   DFF_X1 \buffer_reg[6][2][3][5]  (.D(\input_filter[2][3] [5]), .CK(n_55_6), 
      .Q(\buffer[6][2][3] [5]), .QN());
   DFF_X1 \buffer_reg[6][2][3][4]  (.D(\input_filter[2][3] [4]), .CK(n_55_6), 
      .Q(\buffer[6][2][3] [4]), .QN());
   DFF_X1 \buffer_reg[6][2][3][3]  (.D(\input_filter[2][3] [3]), .CK(n_55_6), 
      .Q(\buffer[6][2][3] [3]), .QN());
   DFF_X1 \buffer_reg[6][2][3][2]  (.D(\input_filter[2][3] [2]), .CK(n_55_6), 
      .Q(\buffer[6][2][3] [2]), .QN());
   DFF_X1 \buffer_reg[6][2][3][1]  (.D(\input_filter[2][3] [1]), .CK(n_55_6), 
      .Q(\buffer[6][2][3] [1]), .QN());
   DFF_X1 \buffer_reg[6][2][3][0]  (.D(\input_filter[2][3] [0]), .CK(n_55_6), 
      .Q(\buffer[6][2][3] [0]), .QN());
   DFF_X1 \buffer_reg[5][2][3][15]  (.D(\input_filter[2][3] [15]), .CK(n_55_7), 
      .Q(\buffer[5][2][3] [15]), .QN());
   DFF_X1 \buffer_reg[5][2][3][14]  (.D(\input_filter[2][3] [14]), .CK(n_55_7), 
      .Q(\buffer[5][2][3] [14]), .QN());
   DFF_X1 \buffer_reg[5][2][3][13]  (.D(\input_filter[2][3] [13]), .CK(n_55_7), 
      .Q(\buffer[5][2][3] [13]), .QN());
   DFF_X1 \buffer_reg[5][2][3][12]  (.D(\input_filter[2][3] [12]), .CK(n_55_7), 
      .Q(\buffer[5][2][3] [12]), .QN());
   DFF_X1 \buffer_reg[5][2][3][11]  (.D(\input_filter[2][3] [11]), .CK(n_55_7), 
      .Q(\buffer[5][2][3] [11]), .QN());
   DFF_X1 \buffer_reg[5][2][3][10]  (.D(\input_filter[2][3] [10]), .CK(n_55_7), 
      .Q(\buffer[5][2][3] [10]), .QN());
   DFF_X1 \buffer_reg[5][2][3][9]  (.D(\input_filter[2][3] [9]), .CK(n_55_7), 
      .Q(\buffer[5][2][3] [9]), .QN());
   DFF_X1 \buffer_reg[5][2][3][8]  (.D(\input_filter[2][3] [8]), .CK(n_55_7), 
      .Q(\buffer[5][2][3] [8]), .QN());
   DFF_X1 \buffer_reg[5][2][3][7]  (.D(\input_filter[2][3] [7]), .CK(n_55_7), 
      .Q(\buffer[5][2][3] [7]), .QN());
   DFF_X1 \buffer_reg[5][2][3][6]  (.D(\input_filter[2][3] [6]), .CK(n_55_7), 
      .Q(\buffer[5][2][3] [6]), .QN());
   DFF_X1 \buffer_reg[5][2][3][5]  (.D(\input_filter[2][3] [5]), .CK(n_55_7), 
      .Q(\buffer[5][2][3] [5]), .QN());
   DFF_X1 \buffer_reg[5][2][3][4]  (.D(\input_filter[2][3] [4]), .CK(n_55_7), 
      .Q(\buffer[5][2][3] [4]), .QN());
   DFF_X1 \buffer_reg[5][2][3][3]  (.D(\input_filter[2][3] [3]), .CK(n_55_7), 
      .Q(\buffer[5][2][3] [3]), .QN());
   DFF_X1 \buffer_reg[5][2][3][2]  (.D(\input_filter[2][3] [2]), .CK(n_55_7), 
      .Q(\buffer[5][2][3] [2]), .QN());
   DFF_X1 \buffer_reg[5][2][3][1]  (.D(\input_filter[2][3] [1]), .CK(n_55_7), 
      .Q(\buffer[5][2][3] [1]), .QN());
   DFF_X1 \buffer_reg[5][2][3][0]  (.D(\input_filter[2][3] [0]), .CK(n_55_7), 
      .Q(\buffer[5][2][3] [0]), .QN());
   DFF_X1 \buffer_reg[4][2][3][15]  (.D(\input_filter[2][3] [15]), .CK(n_55_8), 
      .Q(\buffer[4][2][3] [15]), .QN());
   DFF_X1 \buffer_reg[4][2][3][14]  (.D(\input_filter[2][3] [14]), .CK(n_55_8), 
      .Q(\buffer[4][2][3] [14]), .QN());
   DFF_X1 \buffer_reg[4][2][3][13]  (.D(\input_filter[2][3] [13]), .CK(n_55_8), 
      .Q(\buffer[4][2][3] [13]), .QN());
   DFF_X1 \buffer_reg[4][2][3][12]  (.D(\input_filter[2][3] [12]), .CK(n_55_8), 
      .Q(\buffer[4][2][3] [12]), .QN());
   DFF_X1 \buffer_reg[4][2][3][11]  (.D(\input_filter[2][3] [11]), .CK(n_55_8), 
      .Q(\buffer[4][2][3] [11]), .QN());
   DFF_X1 \buffer_reg[4][2][3][10]  (.D(\input_filter[2][3] [10]), .CK(n_55_8), 
      .Q(\buffer[4][2][3] [10]), .QN());
   DFF_X1 \buffer_reg[4][2][3][9]  (.D(\input_filter[2][3] [9]), .CK(n_55_8), 
      .Q(\buffer[4][2][3] [9]), .QN());
   DFF_X1 \buffer_reg[4][2][3][8]  (.D(\input_filter[2][3] [8]), .CK(n_55_8), 
      .Q(\buffer[4][2][3] [8]), .QN());
   DFF_X1 \buffer_reg[4][2][3][7]  (.D(\input_filter[2][3] [7]), .CK(n_55_8), 
      .Q(\buffer[4][2][3] [7]), .QN());
   DFF_X1 \buffer_reg[4][2][3][6]  (.D(\input_filter[2][3] [6]), .CK(n_55_8), 
      .Q(\buffer[4][2][3] [6]), .QN());
   DFF_X1 \buffer_reg[4][2][3][5]  (.D(\input_filter[2][3] [5]), .CK(n_55_8), 
      .Q(\buffer[4][2][3] [5]), .QN());
   DFF_X1 \buffer_reg[4][2][3][4]  (.D(\input_filter[2][3] [4]), .CK(n_55_8), 
      .Q(\buffer[4][2][3] [4]), .QN());
   DFF_X1 \buffer_reg[4][2][3][3]  (.D(\input_filter[2][3] [3]), .CK(n_55_8), 
      .Q(\buffer[4][2][3] [3]), .QN());
   DFF_X1 \buffer_reg[4][2][3][2]  (.D(\input_filter[2][3] [2]), .CK(n_55_8), 
      .Q(\buffer[4][2][3] [2]), .QN());
   DFF_X1 \buffer_reg[4][2][3][1]  (.D(\input_filter[2][3] [1]), .CK(n_55_8), 
      .Q(\buffer[4][2][3] [1]), .QN());
   DFF_X1 \buffer_reg[4][2][3][0]  (.D(\input_filter[2][3] [0]), .CK(n_55_8), 
      .Q(\buffer[4][2][3] [0]), .QN());
   DFF_X1 \buffer_reg[3][2][3][15]  (.D(\input_filter[2][3] [15]), .CK(n_55_9), 
      .Q(\buffer[3][2][3] [15]), .QN());
   DFF_X1 \buffer_reg[3][2][3][14]  (.D(\input_filter[2][3] [14]), .CK(n_55_9), 
      .Q(\buffer[3][2][3] [14]), .QN());
   DFF_X1 \buffer_reg[3][2][3][13]  (.D(\input_filter[2][3] [13]), .CK(n_55_9), 
      .Q(\buffer[3][2][3] [13]), .QN());
   DFF_X1 \buffer_reg[3][2][3][12]  (.D(\input_filter[2][3] [12]), .CK(n_55_9), 
      .Q(\buffer[3][2][3] [12]), .QN());
   DFF_X1 \buffer_reg[3][2][3][11]  (.D(\input_filter[2][3] [11]), .CK(n_55_9), 
      .Q(\buffer[3][2][3] [11]), .QN());
   DFF_X1 \buffer_reg[3][2][3][10]  (.D(\input_filter[2][3] [10]), .CK(n_55_9), 
      .Q(\buffer[3][2][3] [10]), .QN());
   DFF_X1 \buffer_reg[3][2][3][9]  (.D(\input_filter[2][3] [9]), .CK(n_55_9), 
      .Q(\buffer[3][2][3] [9]), .QN());
   DFF_X1 \buffer_reg[3][2][3][8]  (.D(\input_filter[2][3] [8]), .CK(n_55_9), 
      .Q(\buffer[3][2][3] [8]), .QN());
   DFF_X1 \buffer_reg[3][2][3][7]  (.D(\input_filter[2][3] [7]), .CK(n_55_9), 
      .Q(\buffer[3][2][3] [7]), .QN());
   DFF_X1 \buffer_reg[3][2][3][6]  (.D(\input_filter[2][3] [6]), .CK(n_55_9), 
      .Q(\buffer[3][2][3] [6]), .QN());
   DFF_X1 \buffer_reg[3][2][3][5]  (.D(\input_filter[2][3] [5]), .CK(n_55_9), 
      .Q(\buffer[3][2][3] [5]), .QN());
   DFF_X1 \buffer_reg[3][2][3][4]  (.D(\input_filter[2][3] [4]), .CK(n_55_9), 
      .Q(\buffer[3][2][3] [4]), .QN());
   DFF_X1 \buffer_reg[3][2][3][3]  (.D(\input_filter[2][3] [3]), .CK(n_55_9), 
      .Q(\buffer[3][2][3] [3]), .QN());
   DFF_X1 \buffer_reg[3][2][3][2]  (.D(\input_filter[2][3] [2]), .CK(n_55_9), 
      .Q(\buffer[3][2][3] [2]), .QN());
   DFF_X1 \buffer_reg[3][2][3][1]  (.D(\input_filter[2][3] [1]), .CK(n_55_9), 
      .Q(\buffer[3][2][3] [1]), .QN());
   DFF_X1 \buffer_reg[3][2][3][0]  (.D(\input_filter[2][3] [0]), .CK(n_55_9), 
      .Q(\buffer[3][2][3] [0]), .QN());
   DFF_X1 \buffer_reg[2][2][3][15]  (.D(\input_filter[2][3] [15]), .CK(n_55_10), 
      .Q(\buffer[2][2][3] [15]), .QN());
   DFF_X1 \buffer_reg[2][2][3][14]  (.D(\input_filter[2][3] [14]), .CK(n_55_10), 
      .Q(\buffer[2][2][3] [14]), .QN());
   DFF_X1 \buffer_reg[2][2][3][13]  (.D(\input_filter[2][3] [13]), .CK(n_55_10), 
      .Q(\buffer[2][2][3] [13]), .QN());
   DFF_X1 \buffer_reg[2][2][3][12]  (.D(\input_filter[2][3] [12]), .CK(n_55_10), 
      .Q(\buffer[2][2][3] [12]), .QN());
   DFF_X1 \buffer_reg[2][2][3][11]  (.D(\input_filter[2][3] [11]), .CK(n_55_10), 
      .Q(\buffer[2][2][3] [11]), .QN());
   DFF_X1 \buffer_reg[2][2][3][10]  (.D(\input_filter[2][3] [10]), .CK(n_55_10), 
      .Q(\buffer[2][2][3] [10]), .QN());
   DFF_X1 \buffer_reg[2][2][3][9]  (.D(\input_filter[2][3] [9]), .CK(n_55_10), 
      .Q(\buffer[2][2][3] [9]), .QN());
   DFF_X1 \buffer_reg[2][2][3][8]  (.D(\input_filter[2][3] [8]), .CK(n_55_10), 
      .Q(\buffer[2][2][3] [8]), .QN());
   DFF_X1 \buffer_reg[2][2][3][7]  (.D(\input_filter[2][3] [7]), .CK(n_55_10), 
      .Q(\buffer[2][2][3] [7]), .QN());
   DFF_X1 \buffer_reg[2][2][3][6]  (.D(\input_filter[2][3] [6]), .CK(n_55_10), 
      .Q(\buffer[2][2][3] [6]), .QN());
   DFF_X1 \buffer_reg[2][2][3][5]  (.D(\input_filter[2][3] [5]), .CK(n_55_10), 
      .Q(\buffer[2][2][3] [5]), .QN());
   DFF_X1 \buffer_reg[2][2][3][4]  (.D(\input_filter[2][3] [4]), .CK(n_55_10), 
      .Q(\buffer[2][2][3] [4]), .QN());
   DFF_X1 \buffer_reg[2][2][3][3]  (.D(\input_filter[2][3] [3]), .CK(n_55_10), 
      .Q(\buffer[2][2][3] [3]), .QN());
   DFF_X1 \buffer_reg[2][2][3][2]  (.D(\input_filter[2][3] [2]), .CK(n_55_10), 
      .Q(\buffer[2][2][3] [2]), .QN());
   DFF_X1 \buffer_reg[2][2][3][1]  (.D(\input_filter[2][3] [1]), .CK(n_55_10), 
      .Q(\buffer[2][2][3] [1]), .QN());
   DFF_X1 \buffer_reg[2][2][3][0]  (.D(\input_filter[2][3] [0]), .CK(n_55_10), 
      .Q(\buffer[2][2][3] [0]), .QN());
   DFF_X1 \buffer_reg[1][2][3][15]  (.D(\input_filter[2][3] [15]), .CK(n_55_11), 
      .Q(\buffer[1][2][3] [15]), .QN());
   DFF_X1 \buffer_reg[1][2][3][14]  (.D(\input_filter[2][3] [14]), .CK(n_55_11), 
      .Q(\buffer[1][2][3] [14]), .QN());
   DFF_X1 \buffer_reg[1][2][3][13]  (.D(\input_filter[2][3] [13]), .CK(n_55_11), 
      .Q(\buffer[1][2][3] [13]), .QN());
   DFF_X1 \buffer_reg[1][2][3][12]  (.D(\input_filter[2][3] [12]), .CK(n_55_11), 
      .Q(\buffer[1][2][3] [12]), .QN());
   DFF_X1 \buffer_reg[1][2][3][11]  (.D(\input_filter[2][3] [11]), .CK(n_55_11), 
      .Q(\buffer[1][2][3] [11]), .QN());
   DFF_X1 \buffer_reg[1][2][3][10]  (.D(\input_filter[2][3] [10]), .CK(n_55_11), 
      .Q(\buffer[1][2][3] [10]), .QN());
   DFF_X1 \buffer_reg[1][2][3][9]  (.D(\input_filter[2][3] [9]), .CK(n_55_11), 
      .Q(\buffer[1][2][3] [9]), .QN());
   DFF_X1 \buffer_reg[1][2][3][8]  (.D(\input_filter[2][3] [8]), .CK(n_55_11), 
      .Q(\buffer[1][2][3] [8]), .QN());
   DFF_X1 \buffer_reg[1][2][3][7]  (.D(\input_filter[2][3] [7]), .CK(n_55_11), 
      .Q(\buffer[1][2][3] [7]), .QN());
   DFF_X1 \buffer_reg[1][2][3][6]  (.D(\input_filter[2][3] [6]), .CK(n_55_11), 
      .Q(\buffer[1][2][3] [6]), .QN());
   DFF_X1 \buffer_reg[1][2][3][5]  (.D(\input_filter[2][3] [5]), .CK(n_55_11), 
      .Q(\buffer[1][2][3] [5]), .QN());
   DFF_X1 \buffer_reg[1][2][3][4]  (.D(\input_filter[2][3] [4]), .CK(n_55_11), 
      .Q(\buffer[1][2][3] [4]), .QN());
   DFF_X1 \buffer_reg[1][2][3][3]  (.D(\input_filter[2][3] [3]), .CK(n_55_11), 
      .Q(\buffer[1][2][3] [3]), .QN());
   DFF_X1 \buffer_reg[1][2][3][2]  (.D(\input_filter[2][3] [2]), .CK(n_55_11), 
      .Q(\buffer[1][2][3] [2]), .QN());
   DFF_X1 \buffer_reg[1][2][3][1]  (.D(\input_filter[2][3] [1]), .CK(n_55_11), 
      .Q(\buffer[1][2][3] [1]), .QN());
   DFF_X1 \buffer_reg[1][2][3][0]  (.D(\input_filter[2][3] [0]), .CK(n_55_11), 
      .Q(\buffer[1][2][3] [0]), .QN());
   DFF_X1 \buffer_reg[0][2][3][15]  (.D(\input_filter[2][3] [15]), .CK(n_55_12), 
      .Q(\buffer[0][2][3] [15]), .QN());
   DFF_X1 \buffer_reg[0][2][3][14]  (.D(\input_filter[2][3] [14]), .CK(n_55_12), 
      .Q(\buffer[0][2][3] [14]), .QN());
   DFF_X1 \buffer_reg[0][2][3][13]  (.D(\input_filter[2][3] [13]), .CK(n_55_12), 
      .Q(\buffer[0][2][3] [13]), .QN());
   DFF_X1 \buffer_reg[0][2][3][12]  (.D(\input_filter[2][3] [12]), .CK(n_55_12), 
      .Q(\buffer[0][2][3] [12]), .QN());
   DFF_X1 \buffer_reg[0][2][3][11]  (.D(\input_filter[2][3] [11]), .CK(n_55_12), 
      .Q(\buffer[0][2][3] [11]), .QN());
   DFF_X1 \buffer_reg[0][2][3][10]  (.D(\input_filter[2][3] [10]), .CK(n_55_12), 
      .Q(\buffer[0][2][3] [10]), .QN());
   DFF_X1 \buffer_reg[0][2][3][9]  (.D(\input_filter[2][3] [9]), .CK(n_55_12), 
      .Q(\buffer[0][2][3] [9]), .QN());
   DFF_X1 \buffer_reg[0][2][3][8]  (.D(\input_filter[2][3] [8]), .CK(n_55_12), 
      .Q(\buffer[0][2][3] [8]), .QN());
   DFF_X1 \buffer_reg[0][2][3][7]  (.D(\input_filter[2][3] [7]), .CK(n_55_12), 
      .Q(\buffer[0][2][3] [7]), .QN());
   DFF_X1 \buffer_reg[0][2][3][6]  (.D(\input_filter[2][3] [6]), .CK(n_55_12), 
      .Q(\buffer[0][2][3] [6]), .QN());
   DFF_X1 \buffer_reg[0][2][3][5]  (.D(\input_filter[2][3] [5]), .CK(n_55_12), 
      .Q(\buffer[0][2][3] [5]), .QN());
   DFF_X1 \buffer_reg[0][2][3][4]  (.D(\input_filter[2][3] [4]), .CK(n_55_12), 
      .Q(\buffer[0][2][3] [4]), .QN());
   DFF_X1 \buffer_reg[0][2][3][3]  (.D(\input_filter[2][3] [3]), .CK(n_55_12), 
      .Q(\buffer[0][2][3] [3]), .QN());
   DFF_X1 \buffer_reg[0][2][3][2]  (.D(\input_filter[2][3] [2]), .CK(n_55_12), 
      .Q(\buffer[0][2][3] [2]), .QN());
   DFF_X1 \buffer_reg[0][2][3][1]  (.D(\input_filter[2][3] [1]), .CK(n_55_12), 
      .Q(\buffer[0][2][3] [1]), .QN());
   DFF_X1 \buffer_reg[0][2][3][0]  (.D(\input_filter[2][3] [0]), .CK(n_55_12), 
      .Q(\buffer[0][2][3] [0]), .QN());
   DFF_X1 \buffer_reg[15][2][2][15]  (.D(\input_filter[2][2] [15]), .CK(n_55_13), 
      .Q(\buffer[15][2][2] [15]), .QN());
   DFF_X1 \buffer_reg[15][2][2][14]  (.D(\input_filter[2][2] [14]), .CK(n_55_13), 
      .Q(\buffer[15][2][2] [14]), .QN());
   DFF_X1 \buffer_reg[15][2][2][13]  (.D(\input_filter[2][2] [13]), .CK(n_55_13), 
      .Q(\buffer[15][2][2] [13]), .QN());
   DFF_X1 \buffer_reg[15][2][2][12]  (.D(\input_filter[2][2] [12]), .CK(n_55_13), 
      .Q(\buffer[15][2][2] [12]), .QN());
   DFF_X1 \buffer_reg[15][2][2][11]  (.D(\input_filter[2][2] [11]), .CK(n_55_13), 
      .Q(\buffer[15][2][2] [11]), .QN());
   DFF_X1 \buffer_reg[15][2][2][10]  (.D(\input_filter[2][2] [10]), .CK(n_55_13), 
      .Q(\buffer[15][2][2] [10]), .QN());
   DFF_X1 \buffer_reg[15][2][2][9]  (.D(\input_filter[2][2] [9]), .CK(n_55_13), 
      .Q(\buffer[15][2][2] [9]), .QN());
   DFF_X1 \buffer_reg[15][2][2][8]  (.D(\input_filter[2][2] [8]), .CK(n_55_13), 
      .Q(\buffer[15][2][2] [8]), .QN());
   DFF_X1 \buffer_reg[15][2][2][7]  (.D(\input_filter[2][2] [7]), .CK(n_55_13), 
      .Q(\buffer[15][2][2] [7]), .QN());
   DFF_X1 \buffer_reg[15][2][2][6]  (.D(\input_filter[2][2] [6]), .CK(n_55_13), 
      .Q(\buffer[15][2][2] [6]), .QN());
   DFF_X1 \buffer_reg[15][2][2][5]  (.D(\input_filter[2][2] [5]), .CK(n_55_13), 
      .Q(\buffer[15][2][2] [5]), .QN());
   DFF_X1 \buffer_reg[15][2][2][4]  (.D(\input_filter[2][2] [4]), .CK(n_55_13), 
      .Q(\buffer[15][2][2] [4]), .QN());
   DFF_X1 \buffer_reg[15][2][2][3]  (.D(\input_filter[2][2] [3]), .CK(n_55_13), 
      .Q(\buffer[15][2][2] [3]), .QN());
   DFF_X1 \buffer_reg[15][2][2][2]  (.D(\input_filter[2][2] [2]), .CK(n_55_13), 
      .Q(\buffer[15][2][2] [2]), .QN());
   DFF_X1 \buffer_reg[15][2][2][1]  (.D(\input_filter[2][2] [1]), .CK(n_55_13), 
      .Q(\buffer[15][2][2] [1]), .QN());
   DFF_X1 \buffer_reg[15][2][2][0]  (.D(\input_filter[2][2] [0]), .CK(n_55_13), 
      .Q(\buffer[15][2][2] [0]), .QN());
   DFF_X1 \buffer_reg[14][2][2][15]  (.D(\input_filter[2][2] [15]), .CK(n_55_14), 
      .Q(\buffer[14][2][2] [15]), .QN());
   DFF_X1 \buffer_reg[14][2][2][14]  (.D(\input_filter[2][2] [14]), .CK(n_55_14), 
      .Q(\buffer[14][2][2] [14]), .QN());
   DFF_X1 \buffer_reg[14][2][2][13]  (.D(\input_filter[2][2] [13]), .CK(n_55_14), 
      .Q(\buffer[14][2][2] [13]), .QN());
   DFF_X1 \buffer_reg[14][2][2][12]  (.D(\input_filter[2][2] [12]), .CK(n_55_14), 
      .Q(\buffer[14][2][2] [12]), .QN());
   DFF_X1 \buffer_reg[14][2][2][11]  (.D(\input_filter[2][2] [11]), .CK(n_55_14), 
      .Q(\buffer[14][2][2] [11]), .QN());
   DFF_X1 \buffer_reg[14][2][2][10]  (.D(\input_filter[2][2] [10]), .CK(n_55_14), 
      .Q(\buffer[14][2][2] [10]), .QN());
   DFF_X1 \buffer_reg[14][2][2][9]  (.D(\input_filter[2][2] [9]), .CK(n_55_14), 
      .Q(\buffer[14][2][2] [9]), .QN());
   DFF_X1 \buffer_reg[14][2][2][8]  (.D(\input_filter[2][2] [8]), .CK(n_55_14), 
      .Q(\buffer[14][2][2] [8]), .QN());
   DFF_X1 \buffer_reg[14][2][2][7]  (.D(\input_filter[2][2] [7]), .CK(n_55_14), 
      .Q(\buffer[14][2][2] [7]), .QN());
   DFF_X1 \buffer_reg[14][2][2][6]  (.D(\input_filter[2][2] [6]), .CK(n_55_14), 
      .Q(\buffer[14][2][2] [6]), .QN());
   DFF_X1 \buffer_reg[14][2][2][5]  (.D(\input_filter[2][2] [5]), .CK(n_55_14), 
      .Q(\buffer[14][2][2] [5]), .QN());
   DFF_X1 \buffer_reg[14][2][2][4]  (.D(\input_filter[2][2] [4]), .CK(n_55_14), 
      .Q(\buffer[14][2][2] [4]), .QN());
   DFF_X1 \buffer_reg[14][2][2][3]  (.D(\input_filter[2][2] [3]), .CK(n_55_14), 
      .Q(\buffer[14][2][2] [3]), .QN());
   DFF_X1 \buffer_reg[14][2][2][2]  (.D(\input_filter[2][2] [2]), .CK(n_55_14), 
      .Q(\buffer[14][2][2] [2]), .QN());
   DFF_X1 \buffer_reg[14][2][2][1]  (.D(\input_filter[2][2] [1]), .CK(n_55_14), 
      .Q(\buffer[14][2][2] [1]), .QN());
   DFF_X1 \buffer_reg[14][2][2][0]  (.D(\input_filter[2][2] [0]), .CK(n_55_14), 
      .Q(\buffer[14][2][2] [0]), .QN());
   DFF_X1 \buffer_reg[13][2][2][15]  (.D(\input_filter[2][2] [15]), .CK(n_55_15), 
      .Q(\buffer[13][2][2] [15]), .QN());
   DFF_X1 \buffer_reg[13][2][2][14]  (.D(\input_filter[2][2] [14]), .CK(n_55_15), 
      .Q(\buffer[13][2][2] [14]), .QN());
   DFF_X1 \buffer_reg[13][2][2][13]  (.D(\input_filter[2][2] [13]), .CK(n_55_15), 
      .Q(\buffer[13][2][2] [13]), .QN());
   DFF_X1 \buffer_reg[13][2][2][12]  (.D(\input_filter[2][2] [12]), .CK(n_55_15), 
      .Q(\buffer[13][2][2] [12]), .QN());
   DFF_X1 \buffer_reg[13][2][2][11]  (.D(\input_filter[2][2] [11]), .CK(n_55_15), 
      .Q(\buffer[13][2][2] [11]), .QN());
   DFF_X1 \buffer_reg[13][2][2][10]  (.D(\input_filter[2][2] [10]), .CK(n_55_15), 
      .Q(\buffer[13][2][2] [10]), .QN());
   DFF_X1 \buffer_reg[13][2][2][9]  (.D(\input_filter[2][2] [9]), .CK(n_55_15), 
      .Q(\buffer[13][2][2] [9]), .QN());
   DFF_X1 \buffer_reg[13][2][2][8]  (.D(\input_filter[2][2] [8]), .CK(n_55_15), 
      .Q(\buffer[13][2][2] [8]), .QN());
   DFF_X1 \buffer_reg[13][2][2][7]  (.D(\input_filter[2][2] [7]), .CK(n_55_15), 
      .Q(\buffer[13][2][2] [7]), .QN());
   DFF_X1 \buffer_reg[13][2][2][6]  (.D(\input_filter[2][2] [6]), .CK(n_55_15), 
      .Q(\buffer[13][2][2] [6]), .QN());
   DFF_X1 \buffer_reg[13][2][2][5]  (.D(\input_filter[2][2] [5]), .CK(n_55_15), 
      .Q(\buffer[13][2][2] [5]), .QN());
   DFF_X1 \buffer_reg[13][2][2][4]  (.D(\input_filter[2][2] [4]), .CK(n_55_15), 
      .Q(\buffer[13][2][2] [4]), .QN());
   DFF_X1 \buffer_reg[13][2][2][3]  (.D(\input_filter[2][2] [3]), .CK(n_55_15), 
      .Q(\buffer[13][2][2] [3]), .QN());
   DFF_X1 \buffer_reg[13][2][2][2]  (.D(\input_filter[2][2] [2]), .CK(n_55_15), 
      .Q(\buffer[13][2][2] [2]), .QN());
   DFF_X1 \buffer_reg[13][2][2][1]  (.D(\input_filter[2][2] [1]), .CK(n_55_15), 
      .Q(\buffer[13][2][2] [1]), .QN());
   DFF_X1 \buffer_reg[13][2][2][0]  (.D(\input_filter[2][2] [0]), .CK(n_55_15), 
      .Q(\buffer[13][2][2] [0]), .QN());
   DFF_X1 \buffer_reg[12][2][2][15]  (.D(\input_filter[2][2] [15]), .CK(n_55_0), 
      .Q(\buffer[12][2][2] [15]), .QN());
   DFF_X1 \buffer_reg[12][2][2][14]  (.D(\input_filter[2][2] [14]), .CK(n_55_0), 
      .Q(\buffer[12][2][2] [14]), .QN());
   DFF_X1 \buffer_reg[12][2][2][13]  (.D(\input_filter[2][2] [13]), .CK(n_55_0), 
      .Q(\buffer[12][2][2] [13]), .QN());
   DFF_X1 \buffer_reg[12][2][2][12]  (.D(\input_filter[2][2] [12]), .CK(n_55_0), 
      .Q(\buffer[12][2][2] [12]), .QN());
   DFF_X1 \buffer_reg[12][2][2][11]  (.D(\input_filter[2][2] [11]), .CK(n_55_0), 
      .Q(\buffer[12][2][2] [11]), .QN());
   DFF_X1 \buffer_reg[12][2][2][10]  (.D(\input_filter[2][2] [10]), .CK(n_55_0), 
      .Q(\buffer[12][2][2] [10]), .QN());
   DFF_X1 \buffer_reg[12][2][2][9]  (.D(\input_filter[2][2] [9]), .CK(n_55_0), 
      .Q(\buffer[12][2][2] [9]), .QN());
   DFF_X1 \buffer_reg[12][2][2][8]  (.D(\input_filter[2][2] [8]), .CK(n_55_0), 
      .Q(\buffer[12][2][2] [8]), .QN());
   DFF_X1 \buffer_reg[12][2][2][7]  (.D(\input_filter[2][2] [7]), .CK(n_55_0), 
      .Q(\buffer[12][2][2] [7]), .QN());
   DFF_X1 \buffer_reg[12][2][2][6]  (.D(\input_filter[2][2] [6]), .CK(n_55_0), 
      .Q(\buffer[12][2][2] [6]), .QN());
   DFF_X1 \buffer_reg[12][2][2][5]  (.D(\input_filter[2][2] [5]), .CK(n_55_0), 
      .Q(\buffer[12][2][2] [5]), .QN());
   DFF_X1 \buffer_reg[12][2][2][4]  (.D(\input_filter[2][2] [4]), .CK(n_55_0), 
      .Q(\buffer[12][2][2] [4]), .QN());
   DFF_X1 \buffer_reg[12][2][2][3]  (.D(\input_filter[2][2] [3]), .CK(n_55_0), 
      .Q(\buffer[12][2][2] [3]), .QN());
   DFF_X1 \buffer_reg[12][2][2][2]  (.D(\input_filter[2][2] [2]), .CK(n_55_0), 
      .Q(\buffer[12][2][2] [2]), .QN());
   DFF_X1 \buffer_reg[12][2][2][1]  (.D(\input_filter[2][2] [1]), .CK(n_55_0), 
      .Q(\buffer[12][2][2] [1]), .QN());
   DFF_X1 \buffer_reg[12][2][2][0]  (.D(\input_filter[2][2] [0]), .CK(n_55_0), 
      .Q(\buffer[12][2][2] [0]), .QN());
   DFF_X1 \buffer_reg[11][2][2][15]  (.D(\input_filter[2][2] [15]), .CK(n_55_1), 
      .Q(\buffer[11][2][2] [15]), .QN());
   DFF_X1 \buffer_reg[11][2][2][14]  (.D(\input_filter[2][2] [14]), .CK(n_55_1), 
      .Q(\buffer[11][2][2] [14]), .QN());
   DFF_X1 \buffer_reg[11][2][2][13]  (.D(\input_filter[2][2] [13]), .CK(n_55_1), 
      .Q(\buffer[11][2][2] [13]), .QN());
   DFF_X1 \buffer_reg[11][2][2][12]  (.D(\input_filter[2][2] [12]), .CK(n_55_1), 
      .Q(\buffer[11][2][2] [12]), .QN());
   DFF_X1 \buffer_reg[11][2][2][11]  (.D(\input_filter[2][2] [11]), .CK(n_55_1), 
      .Q(\buffer[11][2][2] [11]), .QN());
   DFF_X1 \buffer_reg[11][2][2][10]  (.D(\input_filter[2][2] [10]), .CK(n_55_1), 
      .Q(\buffer[11][2][2] [10]), .QN());
   DFF_X1 \buffer_reg[11][2][2][9]  (.D(\input_filter[2][2] [9]), .CK(n_55_1), 
      .Q(\buffer[11][2][2] [9]), .QN());
   DFF_X1 \buffer_reg[11][2][2][8]  (.D(\input_filter[2][2] [8]), .CK(n_55_1), 
      .Q(\buffer[11][2][2] [8]), .QN());
   DFF_X1 \buffer_reg[11][2][2][7]  (.D(\input_filter[2][2] [7]), .CK(n_55_1), 
      .Q(\buffer[11][2][2] [7]), .QN());
   DFF_X1 \buffer_reg[11][2][2][6]  (.D(\input_filter[2][2] [6]), .CK(n_55_1), 
      .Q(\buffer[11][2][2] [6]), .QN());
   DFF_X1 \buffer_reg[11][2][2][5]  (.D(\input_filter[2][2] [5]), .CK(n_55_1), 
      .Q(\buffer[11][2][2] [5]), .QN());
   DFF_X1 \buffer_reg[11][2][2][4]  (.D(\input_filter[2][2] [4]), .CK(n_55_1), 
      .Q(\buffer[11][2][2] [4]), .QN());
   DFF_X1 \buffer_reg[11][2][2][3]  (.D(\input_filter[2][2] [3]), .CK(n_55_1), 
      .Q(\buffer[11][2][2] [3]), .QN());
   DFF_X1 \buffer_reg[11][2][2][2]  (.D(\input_filter[2][2] [2]), .CK(n_55_1), 
      .Q(\buffer[11][2][2] [2]), .QN());
   DFF_X1 \buffer_reg[11][2][2][1]  (.D(\input_filter[2][2] [1]), .CK(n_55_1), 
      .Q(\buffer[11][2][2] [1]), .QN());
   DFF_X1 \buffer_reg[11][2][2][0]  (.D(\input_filter[2][2] [0]), .CK(n_55_1), 
      .Q(\buffer[11][2][2] [0]), .QN());
   DFF_X1 \buffer_reg[10][2][2][15]  (.D(\input_filter[2][2] [15]), .CK(n_55_2), 
      .Q(\buffer[10][2][2] [15]), .QN());
   DFF_X1 \buffer_reg[10][2][2][14]  (.D(\input_filter[2][2] [14]), .CK(n_55_2), 
      .Q(\buffer[10][2][2] [14]), .QN());
   DFF_X1 \buffer_reg[10][2][2][13]  (.D(\input_filter[2][2] [13]), .CK(n_55_2), 
      .Q(\buffer[10][2][2] [13]), .QN());
   DFF_X1 \buffer_reg[10][2][2][12]  (.D(\input_filter[2][2] [12]), .CK(n_55_2), 
      .Q(\buffer[10][2][2] [12]), .QN());
   DFF_X1 \buffer_reg[10][2][2][11]  (.D(\input_filter[2][2] [11]), .CK(n_55_2), 
      .Q(\buffer[10][2][2] [11]), .QN());
   DFF_X1 \buffer_reg[10][2][2][10]  (.D(\input_filter[2][2] [10]), .CK(n_55_2), 
      .Q(\buffer[10][2][2] [10]), .QN());
   DFF_X1 \buffer_reg[10][2][2][9]  (.D(\input_filter[2][2] [9]), .CK(n_55_2), 
      .Q(\buffer[10][2][2] [9]), .QN());
   DFF_X1 \buffer_reg[10][2][2][8]  (.D(\input_filter[2][2] [8]), .CK(n_55_2), 
      .Q(\buffer[10][2][2] [8]), .QN());
   DFF_X1 \buffer_reg[10][2][2][7]  (.D(\input_filter[2][2] [7]), .CK(n_55_2), 
      .Q(\buffer[10][2][2] [7]), .QN());
   DFF_X1 \buffer_reg[10][2][2][6]  (.D(\input_filter[2][2] [6]), .CK(n_55_2), 
      .Q(\buffer[10][2][2] [6]), .QN());
   DFF_X1 \buffer_reg[10][2][2][5]  (.D(\input_filter[2][2] [5]), .CK(n_55_2), 
      .Q(\buffer[10][2][2] [5]), .QN());
   DFF_X1 \buffer_reg[10][2][2][4]  (.D(\input_filter[2][2] [4]), .CK(n_55_2), 
      .Q(\buffer[10][2][2] [4]), .QN());
   DFF_X1 \buffer_reg[10][2][2][3]  (.D(\input_filter[2][2] [3]), .CK(n_55_2), 
      .Q(\buffer[10][2][2] [3]), .QN());
   DFF_X1 \buffer_reg[10][2][2][2]  (.D(\input_filter[2][2] [2]), .CK(n_55_2), 
      .Q(\buffer[10][2][2] [2]), .QN());
   DFF_X1 \buffer_reg[10][2][2][1]  (.D(\input_filter[2][2] [1]), .CK(n_55_2), 
      .Q(\buffer[10][2][2] [1]), .QN());
   DFF_X1 \buffer_reg[10][2][2][0]  (.D(\input_filter[2][2] [0]), .CK(n_55_2), 
      .Q(\buffer[10][2][2] [0]), .QN());
   DFF_X1 \buffer_reg[9][2][2][15]  (.D(\input_filter[2][2] [15]), .CK(n_55_3), 
      .Q(\buffer[9][2][2] [15]), .QN());
   DFF_X1 \buffer_reg[9][2][2][14]  (.D(\input_filter[2][2] [14]), .CK(n_55_3), 
      .Q(\buffer[9][2][2] [14]), .QN());
   DFF_X1 \buffer_reg[9][2][2][13]  (.D(\input_filter[2][2] [13]), .CK(n_55_3), 
      .Q(\buffer[9][2][2] [13]), .QN());
   DFF_X1 \buffer_reg[9][2][2][12]  (.D(\input_filter[2][2] [12]), .CK(n_55_3), 
      .Q(\buffer[9][2][2] [12]), .QN());
   DFF_X1 \buffer_reg[9][2][2][11]  (.D(\input_filter[2][2] [11]), .CK(n_55_3), 
      .Q(\buffer[9][2][2] [11]), .QN());
   DFF_X1 \buffer_reg[9][2][2][10]  (.D(\input_filter[2][2] [10]), .CK(n_55_3), 
      .Q(\buffer[9][2][2] [10]), .QN());
   DFF_X1 \buffer_reg[9][2][2][9]  (.D(\input_filter[2][2] [9]), .CK(n_55_3), 
      .Q(\buffer[9][2][2] [9]), .QN());
   DFF_X1 \buffer_reg[9][2][2][8]  (.D(\input_filter[2][2] [8]), .CK(n_55_3), 
      .Q(\buffer[9][2][2] [8]), .QN());
   DFF_X1 \buffer_reg[9][2][2][7]  (.D(\input_filter[2][2] [7]), .CK(n_55_3), 
      .Q(\buffer[9][2][2] [7]), .QN());
   DFF_X1 \buffer_reg[9][2][2][6]  (.D(\input_filter[2][2] [6]), .CK(n_55_3), 
      .Q(\buffer[9][2][2] [6]), .QN());
   DFF_X1 \buffer_reg[9][2][2][5]  (.D(\input_filter[2][2] [5]), .CK(n_55_3), 
      .Q(\buffer[9][2][2] [5]), .QN());
   DFF_X1 \buffer_reg[9][2][2][4]  (.D(\input_filter[2][2] [4]), .CK(n_55_3), 
      .Q(\buffer[9][2][2] [4]), .QN());
   DFF_X1 \buffer_reg[9][2][2][3]  (.D(\input_filter[2][2] [3]), .CK(n_55_3), 
      .Q(\buffer[9][2][2] [3]), .QN());
   DFF_X1 \buffer_reg[9][2][2][2]  (.D(\input_filter[2][2] [2]), .CK(n_55_3), 
      .Q(\buffer[9][2][2] [2]), .QN());
   DFF_X1 \buffer_reg[9][2][2][1]  (.D(\input_filter[2][2] [1]), .CK(n_55_3), 
      .Q(\buffer[9][2][2] [1]), .QN());
   DFF_X1 \buffer_reg[9][2][2][0]  (.D(\input_filter[2][2] [0]), .CK(n_55_3), 
      .Q(\buffer[9][2][2] [0]), .QN());
   DFF_X1 \buffer_reg[8][2][2][15]  (.D(\input_filter[2][2] [15]), .CK(n_55_4), 
      .Q(\buffer[8][2][2] [15]), .QN());
   DFF_X1 \buffer_reg[8][2][2][14]  (.D(\input_filter[2][2] [14]), .CK(n_55_4), 
      .Q(\buffer[8][2][2] [14]), .QN());
   DFF_X1 \buffer_reg[8][2][2][13]  (.D(\input_filter[2][2] [13]), .CK(n_55_4), 
      .Q(\buffer[8][2][2] [13]), .QN());
   DFF_X1 \buffer_reg[8][2][2][12]  (.D(\input_filter[2][2] [12]), .CK(n_55_4), 
      .Q(\buffer[8][2][2] [12]), .QN());
   DFF_X1 \buffer_reg[8][2][2][11]  (.D(\input_filter[2][2] [11]), .CK(n_55_4), 
      .Q(\buffer[8][2][2] [11]), .QN());
   DFF_X1 \buffer_reg[8][2][2][10]  (.D(\input_filter[2][2] [10]), .CK(n_55_4), 
      .Q(\buffer[8][2][2] [10]), .QN());
   DFF_X1 \buffer_reg[8][2][2][9]  (.D(\input_filter[2][2] [9]), .CK(n_55_4), 
      .Q(\buffer[8][2][2] [9]), .QN());
   DFF_X1 \buffer_reg[8][2][2][8]  (.D(\input_filter[2][2] [8]), .CK(n_55_4), 
      .Q(\buffer[8][2][2] [8]), .QN());
   DFF_X1 \buffer_reg[8][2][2][7]  (.D(\input_filter[2][2] [7]), .CK(n_55_4), 
      .Q(\buffer[8][2][2] [7]), .QN());
   DFF_X1 \buffer_reg[8][2][2][6]  (.D(\input_filter[2][2] [6]), .CK(n_55_4), 
      .Q(\buffer[8][2][2] [6]), .QN());
   DFF_X1 \buffer_reg[8][2][2][5]  (.D(\input_filter[2][2] [5]), .CK(n_55_4), 
      .Q(\buffer[8][2][2] [5]), .QN());
   DFF_X1 \buffer_reg[8][2][2][4]  (.D(\input_filter[2][2] [4]), .CK(n_55_4), 
      .Q(\buffer[8][2][2] [4]), .QN());
   DFF_X1 \buffer_reg[8][2][2][3]  (.D(\input_filter[2][2] [3]), .CK(n_55_4), 
      .Q(\buffer[8][2][2] [3]), .QN());
   DFF_X1 \buffer_reg[8][2][2][2]  (.D(\input_filter[2][2] [2]), .CK(n_55_4), 
      .Q(\buffer[8][2][2] [2]), .QN());
   DFF_X1 \buffer_reg[8][2][2][1]  (.D(\input_filter[2][2] [1]), .CK(n_55_4), 
      .Q(\buffer[8][2][2] [1]), .QN());
   DFF_X1 \buffer_reg[8][2][2][0]  (.D(\input_filter[2][2] [0]), .CK(n_55_4), 
      .Q(\buffer[8][2][2] [0]), .QN());
   DFF_X1 \buffer_reg[7][2][2][15]  (.D(\input_filter[2][2] [15]), .CK(n_55_5), 
      .Q(\buffer[7][2][2] [15]), .QN());
   DFF_X1 \buffer_reg[7][2][2][14]  (.D(\input_filter[2][2] [14]), .CK(n_55_5), 
      .Q(\buffer[7][2][2] [14]), .QN());
   DFF_X1 \buffer_reg[7][2][2][13]  (.D(\input_filter[2][2] [13]), .CK(n_55_5), 
      .Q(\buffer[7][2][2] [13]), .QN());
   DFF_X1 \buffer_reg[7][2][2][12]  (.D(\input_filter[2][2] [12]), .CK(n_55_5), 
      .Q(\buffer[7][2][2] [12]), .QN());
   DFF_X1 \buffer_reg[7][2][2][11]  (.D(\input_filter[2][2] [11]), .CK(n_55_5), 
      .Q(\buffer[7][2][2] [11]), .QN());
   DFF_X1 \buffer_reg[7][2][2][10]  (.D(\input_filter[2][2] [10]), .CK(n_55_5), 
      .Q(\buffer[7][2][2] [10]), .QN());
   DFF_X1 \buffer_reg[7][2][2][9]  (.D(\input_filter[2][2] [9]), .CK(n_55_5), 
      .Q(\buffer[7][2][2] [9]), .QN());
   DFF_X1 \buffer_reg[7][2][2][8]  (.D(\input_filter[2][2] [8]), .CK(n_55_5), 
      .Q(\buffer[7][2][2] [8]), .QN());
   DFF_X1 \buffer_reg[7][2][2][7]  (.D(\input_filter[2][2] [7]), .CK(n_55_5), 
      .Q(\buffer[7][2][2] [7]), .QN());
   DFF_X1 \buffer_reg[7][2][2][6]  (.D(\input_filter[2][2] [6]), .CK(n_55_5), 
      .Q(\buffer[7][2][2] [6]), .QN());
   DFF_X1 \buffer_reg[7][2][2][5]  (.D(\input_filter[2][2] [5]), .CK(n_55_5), 
      .Q(\buffer[7][2][2] [5]), .QN());
   DFF_X1 \buffer_reg[7][2][2][4]  (.D(\input_filter[2][2] [4]), .CK(n_55_5), 
      .Q(\buffer[7][2][2] [4]), .QN());
   DFF_X1 \buffer_reg[7][2][2][3]  (.D(\input_filter[2][2] [3]), .CK(n_55_5), 
      .Q(\buffer[7][2][2] [3]), .QN());
   DFF_X1 \buffer_reg[7][2][2][2]  (.D(\input_filter[2][2] [2]), .CK(n_55_5), 
      .Q(\buffer[7][2][2] [2]), .QN());
   DFF_X1 \buffer_reg[7][2][2][1]  (.D(\input_filter[2][2] [1]), .CK(n_55_5), 
      .Q(\buffer[7][2][2] [1]), .QN());
   DFF_X1 \buffer_reg[7][2][2][0]  (.D(\input_filter[2][2] [0]), .CK(n_55_5), 
      .Q(\buffer[7][2][2] [0]), .QN());
   DFF_X1 \buffer_reg[6][2][2][15]  (.D(\input_filter[2][2] [15]), .CK(n_55_6), 
      .Q(\buffer[6][2][2] [15]), .QN());
   DFF_X1 \buffer_reg[6][2][2][14]  (.D(\input_filter[2][2] [14]), .CK(n_55_6), 
      .Q(\buffer[6][2][2] [14]), .QN());
   DFF_X1 \buffer_reg[6][2][2][13]  (.D(\input_filter[2][2] [13]), .CK(n_55_6), 
      .Q(\buffer[6][2][2] [13]), .QN());
   DFF_X1 \buffer_reg[6][2][2][12]  (.D(\input_filter[2][2] [12]), .CK(n_55_6), 
      .Q(\buffer[6][2][2] [12]), .QN());
   DFF_X1 \buffer_reg[6][2][2][11]  (.D(\input_filter[2][2] [11]), .CK(n_55_6), 
      .Q(\buffer[6][2][2] [11]), .QN());
   DFF_X1 \buffer_reg[6][2][2][10]  (.D(\input_filter[2][2] [10]), .CK(n_55_6), 
      .Q(\buffer[6][2][2] [10]), .QN());
   DFF_X1 \buffer_reg[6][2][2][9]  (.D(\input_filter[2][2] [9]), .CK(n_55_6), 
      .Q(\buffer[6][2][2] [9]), .QN());
   DFF_X1 \buffer_reg[6][2][2][8]  (.D(\input_filter[2][2] [8]), .CK(n_55_6), 
      .Q(\buffer[6][2][2] [8]), .QN());
   DFF_X1 \buffer_reg[6][2][2][7]  (.D(\input_filter[2][2] [7]), .CK(n_55_6), 
      .Q(\buffer[6][2][2] [7]), .QN());
   DFF_X1 \buffer_reg[6][2][2][6]  (.D(\input_filter[2][2] [6]), .CK(n_55_6), 
      .Q(\buffer[6][2][2] [6]), .QN());
   DFF_X1 \buffer_reg[6][2][2][5]  (.D(\input_filter[2][2] [5]), .CK(n_55_6), 
      .Q(\buffer[6][2][2] [5]), .QN());
   DFF_X1 \buffer_reg[6][2][2][4]  (.D(\input_filter[2][2] [4]), .CK(n_55_6), 
      .Q(\buffer[6][2][2] [4]), .QN());
   DFF_X1 \buffer_reg[6][2][2][3]  (.D(\input_filter[2][2] [3]), .CK(n_55_6), 
      .Q(\buffer[6][2][2] [3]), .QN());
   DFF_X1 \buffer_reg[6][2][2][2]  (.D(\input_filter[2][2] [2]), .CK(n_55_6), 
      .Q(\buffer[6][2][2] [2]), .QN());
   DFF_X1 \buffer_reg[6][2][2][1]  (.D(\input_filter[2][2] [1]), .CK(n_55_6), 
      .Q(\buffer[6][2][2] [1]), .QN());
   DFF_X1 \buffer_reg[6][2][2][0]  (.D(\input_filter[2][2] [0]), .CK(n_55_6), 
      .Q(\buffer[6][2][2] [0]), .QN());
   DFF_X1 \buffer_reg[5][2][2][15]  (.D(\input_filter[2][2] [15]), .CK(n_55_7), 
      .Q(\buffer[5][2][2] [15]), .QN());
   DFF_X1 \buffer_reg[5][2][2][14]  (.D(\input_filter[2][2] [14]), .CK(n_55_7), 
      .Q(\buffer[5][2][2] [14]), .QN());
   DFF_X1 \buffer_reg[5][2][2][13]  (.D(\input_filter[2][2] [13]), .CK(n_55_7), 
      .Q(\buffer[5][2][2] [13]), .QN());
   DFF_X1 \buffer_reg[5][2][2][12]  (.D(\input_filter[2][2] [12]), .CK(n_55_7), 
      .Q(\buffer[5][2][2] [12]), .QN());
   DFF_X1 \buffer_reg[5][2][2][11]  (.D(\input_filter[2][2] [11]), .CK(n_55_7), 
      .Q(\buffer[5][2][2] [11]), .QN());
   DFF_X1 \buffer_reg[5][2][2][10]  (.D(\input_filter[2][2] [10]), .CK(n_55_7), 
      .Q(\buffer[5][2][2] [10]), .QN());
   DFF_X1 \buffer_reg[5][2][2][9]  (.D(\input_filter[2][2] [9]), .CK(n_55_7), 
      .Q(\buffer[5][2][2] [9]), .QN());
   DFF_X1 \buffer_reg[5][2][2][8]  (.D(\input_filter[2][2] [8]), .CK(n_55_7), 
      .Q(\buffer[5][2][2] [8]), .QN());
   DFF_X1 \buffer_reg[5][2][2][7]  (.D(\input_filter[2][2] [7]), .CK(n_55_7), 
      .Q(\buffer[5][2][2] [7]), .QN());
   DFF_X1 \buffer_reg[5][2][2][6]  (.D(\input_filter[2][2] [6]), .CK(n_55_7), 
      .Q(\buffer[5][2][2] [6]), .QN());
   DFF_X1 \buffer_reg[5][2][2][5]  (.D(\input_filter[2][2] [5]), .CK(n_55_7), 
      .Q(\buffer[5][2][2] [5]), .QN());
   DFF_X1 \buffer_reg[5][2][2][4]  (.D(\input_filter[2][2] [4]), .CK(n_55_7), 
      .Q(\buffer[5][2][2] [4]), .QN());
   DFF_X1 \buffer_reg[5][2][2][3]  (.D(\input_filter[2][2] [3]), .CK(n_55_7), 
      .Q(\buffer[5][2][2] [3]), .QN());
   DFF_X1 \buffer_reg[5][2][2][2]  (.D(\input_filter[2][2] [2]), .CK(n_55_7), 
      .Q(\buffer[5][2][2] [2]), .QN());
   DFF_X1 \buffer_reg[5][2][2][1]  (.D(\input_filter[2][2] [1]), .CK(n_55_7), 
      .Q(\buffer[5][2][2] [1]), .QN());
   DFF_X1 \buffer_reg[5][2][2][0]  (.D(\input_filter[2][2] [0]), .CK(n_55_7), 
      .Q(\buffer[5][2][2] [0]), .QN());
   DFF_X1 \buffer_reg[4][2][2][15]  (.D(\input_filter[2][2] [15]), .CK(n_55_8), 
      .Q(\buffer[4][2][2] [15]), .QN());
   DFF_X1 \buffer_reg[4][2][2][14]  (.D(\input_filter[2][2] [14]), .CK(n_55_8), 
      .Q(\buffer[4][2][2] [14]), .QN());
   DFF_X1 \buffer_reg[4][2][2][13]  (.D(\input_filter[2][2] [13]), .CK(n_55_8), 
      .Q(\buffer[4][2][2] [13]), .QN());
   DFF_X1 \buffer_reg[4][2][2][12]  (.D(\input_filter[2][2] [12]), .CK(n_55_8), 
      .Q(\buffer[4][2][2] [12]), .QN());
   DFF_X1 \buffer_reg[4][2][2][11]  (.D(\input_filter[2][2] [11]), .CK(n_55_8), 
      .Q(\buffer[4][2][2] [11]), .QN());
   DFF_X1 \buffer_reg[4][2][2][10]  (.D(\input_filter[2][2] [10]), .CK(n_55_8), 
      .Q(\buffer[4][2][2] [10]), .QN());
   DFF_X1 \buffer_reg[4][2][2][9]  (.D(\input_filter[2][2] [9]), .CK(n_55_8), 
      .Q(\buffer[4][2][2] [9]), .QN());
   DFF_X1 \buffer_reg[4][2][2][8]  (.D(\input_filter[2][2] [8]), .CK(n_55_8), 
      .Q(\buffer[4][2][2] [8]), .QN());
   DFF_X1 \buffer_reg[4][2][2][7]  (.D(\input_filter[2][2] [7]), .CK(n_55_8), 
      .Q(\buffer[4][2][2] [7]), .QN());
   DFF_X1 \buffer_reg[4][2][2][6]  (.D(\input_filter[2][2] [6]), .CK(n_55_8), 
      .Q(\buffer[4][2][2] [6]), .QN());
   DFF_X1 \buffer_reg[4][2][2][5]  (.D(\input_filter[2][2] [5]), .CK(n_55_8), 
      .Q(\buffer[4][2][2] [5]), .QN());
   DFF_X1 \buffer_reg[4][2][2][4]  (.D(\input_filter[2][2] [4]), .CK(n_55_8), 
      .Q(\buffer[4][2][2] [4]), .QN());
   DFF_X1 \buffer_reg[4][2][2][3]  (.D(\input_filter[2][2] [3]), .CK(n_55_8), 
      .Q(\buffer[4][2][2] [3]), .QN());
   DFF_X1 \buffer_reg[4][2][2][2]  (.D(\input_filter[2][2] [2]), .CK(n_55_8), 
      .Q(\buffer[4][2][2] [2]), .QN());
   DFF_X1 \buffer_reg[4][2][2][1]  (.D(\input_filter[2][2] [1]), .CK(n_55_8), 
      .Q(\buffer[4][2][2] [1]), .QN());
   DFF_X1 \buffer_reg[4][2][2][0]  (.D(\input_filter[2][2] [0]), .CK(n_55_8), 
      .Q(\buffer[4][2][2] [0]), .QN());
   DFF_X1 \buffer_reg[3][2][2][15]  (.D(\input_filter[2][2] [15]), .CK(n_55_9), 
      .Q(\buffer[3][2][2] [15]), .QN());
   DFF_X1 \buffer_reg[3][2][2][14]  (.D(\input_filter[2][2] [14]), .CK(n_55_9), 
      .Q(\buffer[3][2][2] [14]), .QN());
   DFF_X1 \buffer_reg[3][2][2][13]  (.D(\input_filter[2][2] [13]), .CK(n_55_9), 
      .Q(\buffer[3][2][2] [13]), .QN());
   DFF_X1 \buffer_reg[3][2][2][12]  (.D(\input_filter[2][2] [12]), .CK(n_55_9), 
      .Q(\buffer[3][2][2] [12]), .QN());
   DFF_X1 \buffer_reg[3][2][2][11]  (.D(\input_filter[2][2] [11]), .CK(n_55_9), 
      .Q(\buffer[3][2][2] [11]), .QN());
   DFF_X1 \buffer_reg[3][2][2][10]  (.D(\input_filter[2][2] [10]), .CK(n_55_9), 
      .Q(\buffer[3][2][2] [10]), .QN());
   DFF_X1 \buffer_reg[3][2][2][9]  (.D(\input_filter[2][2] [9]), .CK(n_55_9), 
      .Q(\buffer[3][2][2] [9]), .QN());
   DFF_X1 \buffer_reg[3][2][2][8]  (.D(\input_filter[2][2] [8]), .CK(n_55_9), 
      .Q(\buffer[3][2][2] [8]), .QN());
   DFF_X1 \buffer_reg[3][2][2][7]  (.D(\input_filter[2][2] [7]), .CK(n_55_9), 
      .Q(\buffer[3][2][2] [7]), .QN());
   DFF_X1 \buffer_reg[3][2][2][6]  (.D(\input_filter[2][2] [6]), .CK(n_55_9), 
      .Q(\buffer[3][2][2] [6]), .QN());
   DFF_X1 \buffer_reg[3][2][2][5]  (.D(\input_filter[2][2] [5]), .CK(n_55_9), 
      .Q(\buffer[3][2][2] [5]), .QN());
   DFF_X1 \buffer_reg[3][2][2][4]  (.D(\input_filter[2][2] [4]), .CK(n_55_9), 
      .Q(\buffer[3][2][2] [4]), .QN());
   DFF_X1 \buffer_reg[3][2][2][3]  (.D(\input_filter[2][2] [3]), .CK(n_55_9), 
      .Q(\buffer[3][2][2] [3]), .QN());
   DFF_X1 \buffer_reg[3][2][2][2]  (.D(\input_filter[2][2] [2]), .CK(n_55_9), 
      .Q(\buffer[3][2][2] [2]), .QN());
   DFF_X1 \buffer_reg[3][2][2][1]  (.D(\input_filter[2][2] [1]), .CK(n_55_9), 
      .Q(\buffer[3][2][2] [1]), .QN());
   DFF_X1 \buffer_reg[3][2][2][0]  (.D(\input_filter[2][2] [0]), .CK(n_55_9), 
      .Q(\buffer[3][2][2] [0]), .QN());
   DFF_X1 \buffer_reg[2][2][2][15]  (.D(\input_filter[2][2] [15]), .CK(n_55_10), 
      .Q(\buffer[2][2][2] [15]), .QN());
   DFF_X1 \buffer_reg[2][2][2][14]  (.D(\input_filter[2][2] [14]), .CK(n_55_10), 
      .Q(\buffer[2][2][2] [14]), .QN());
   DFF_X1 \buffer_reg[2][2][2][13]  (.D(\input_filter[2][2] [13]), .CK(n_55_10), 
      .Q(\buffer[2][2][2] [13]), .QN());
   DFF_X1 \buffer_reg[2][2][2][12]  (.D(\input_filter[2][2] [12]), .CK(n_55_10), 
      .Q(\buffer[2][2][2] [12]), .QN());
   DFF_X1 \buffer_reg[2][2][2][11]  (.D(\input_filter[2][2] [11]), .CK(n_55_10), 
      .Q(\buffer[2][2][2] [11]), .QN());
   DFF_X1 \buffer_reg[2][2][2][10]  (.D(\input_filter[2][2] [10]), .CK(n_55_10), 
      .Q(\buffer[2][2][2] [10]), .QN());
   DFF_X1 \buffer_reg[2][2][2][9]  (.D(\input_filter[2][2] [9]), .CK(n_55_10), 
      .Q(\buffer[2][2][2] [9]), .QN());
   DFF_X1 \buffer_reg[2][2][2][8]  (.D(\input_filter[2][2] [8]), .CK(n_55_10), 
      .Q(\buffer[2][2][2] [8]), .QN());
   DFF_X1 \buffer_reg[2][2][2][7]  (.D(\input_filter[2][2] [7]), .CK(n_55_10), 
      .Q(\buffer[2][2][2] [7]), .QN());
   DFF_X1 \buffer_reg[2][2][2][6]  (.D(\input_filter[2][2] [6]), .CK(n_55_10), 
      .Q(\buffer[2][2][2] [6]), .QN());
   DFF_X1 \buffer_reg[2][2][2][5]  (.D(\input_filter[2][2] [5]), .CK(n_55_10), 
      .Q(\buffer[2][2][2] [5]), .QN());
   DFF_X1 \buffer_reg[2][2][2][4]  (.D(\input_filter[2][2] [4]), .CK(n_55_10), 
      .Q(\buffer[2][2][2] [4]), .QN());
   DFF_X1 \buffer_reg[2][2][2][3]  (.D(\input_filter[2][2] [3]), .CK(n_55_10), 
      .Q(\buffer[2][2][2] [3]), .QN());
   DFF_X1 \buffer_reg[2][2][2][2]  (.D(\input_filter[2][2] [2]), .CK(n_55_10), 
      .Q(\buffer[2][2][2] [2]), .QN());
   DFF_X1 \buffer_reg[2][2][2][1]  (.D(\input_filter[2][2] [1]), .CK(n_55_10), 
      .Q(\buffer[2][2][2] [1]), .QN());
   DFF_X1 \buffer_reg[2][2][2][0]  (.D(\input_filter[2][2] [0]), .CK(n_55_10), 
      .Q(\buffer[2][2][2] [0]), .QN());
   DFF_X1 \buffer_reg[1][2][2][15]  (.D(\input_filter[2][2] [15]), .CK(n_55_11), 
      .Q(\buffer[1][2][2] [15]), .QN());
   DFF_X1 \buffer_reg[1][2][2][14]  (.D(\input_filter[2][2] [14]), .CK(n_55_11), 
      .Q(\buffer[1][2][2] [14]), .QN());
   DFF_X1 \buffer_reg[1][2][2][13]  (.D(\input_filter[2][2] [13]), .CK(n_55_11), 
      .Q(\buffer[1][2][2] [13]), .QN());
   DFF_X1 \buffer_reg[1][2][2][12]  (.D(\input_filter[2][2] [12]), .CK(n_55_11), 
      .Q(\buffer[1][2][2] [12]), .QN());
   DFF_X1 \buffer_reg[1][2][2][11]  (.D(\input_filter[2][2] [11]), .CK(n_55_11), 
      .Q(\buffer[1][2][2] [11]), .QN());
   DFF_X1 \buffer_reg[1][2][2][10]  (.D(\input_filter[2][2] [10]), .CK(n_55_11), 
      .Q(\buffer[1][2][2] [10]), .QN());
   DFF_X1 \buffer_reg[1][2][2][9]  (.D(\input_filter[2][2] [9]), .CK(n_55_11), 
      .Q(\buffer[1][2][2] [9]), .QN());
   DFF_X1 \buffer_reg[1][2][2][8]  (.D(\input_filter[2][2] [8]), .CK(n_55_11), 
      .Q(\buffer[1][2][2] [8]), .QN());
   DFF_X1 \buffer_reg[1][2][2][7]  (.D(\input_filter[2][2] [7]), .CK(n_55_11), 
      .Q(\buffer[1][2][2] [7]), .QN());
   DFF_X1 \buffer_reg[1][2][2][6]  (.D(\input_filter[2][2] [6]), .CK(n_55_11), 
      .Q(\buffer[1][2][2] [6]), .QN());
   DFF_X1 \buffer_reg[1][2][2][5]  (.D(\input_filter[2][2] [5]), .CK(n_55_11), 
      .Q(\buffer[1][2][2] [5]), .QN());
   DFF_X1 \buffer_reg[1][2][2][4]  (.D(\input_filter[2][2] [4]), .CK(n_55_11), 
      .Q(\buffer[1][2][2] [4]), .QN());
   DFF_X1 \buffer_reg[1][2][2][3]  (.D(\input_filter[2][2] [3]), .CK(n_55_11), 
      .Q(\buffer[1][2][2] [3]), .QN());
   DFF_X1 \buffer_reg[1][2][2][2]  (.D(\input_filter[2][2] [2]), .CK(n_55_11), 
      .Q(\buffer[1][2][2] [2]), .QN());
   DFF_X1 \buffer_reg[1][2][2][1]  (.D(\input_filter[2][2] [1]), .CK(n_55_11), 
      .Q(\buffer[1][2][2] [1]), .QN());
   DFF_X1 \buffer_reg[1][2][2][0]  (.D(\input_filter[2][2] [0]), .CK(n_55_11), 
      .Q(\buffer[1][2][2] [0]), .QN());
   DFF_X1 \buffer_reg[0][2][2][15]  (.D(\input_filter[2][2] [15]), .CK(n_55_12), 
      .Q(\buffer[0][2][2] [15]), .QN());
   DFF_X1 \buffer_reg[0][2][2][14]  (.D(\input_filter[2][2] [14]), .CK(n_55_12), 
      .Q(\buffer[0][2][2] [14]), .QN());
   DFF_X1 \buffer_reg[0][2][2][13]  (.D(\input_filter[2][2] [13]), .CK(n_55_12), 
      .Q(\buffer[0][2][2] [13]), .QN());
   DFF_X1 \buffer_reg[0][2][2][12]  (.D(\input_filter[2][2] [12]), .CK(n_55_12), 
      .Q(\buffer[0][2][2] [12]), .QN());
   DFF_X1 \buffer_reg[0][2][2][11]  (.D(\input_filter[2][2] [11]), .CK(n_55_12), 
      .Q(\buffer[0][2][2] [11]), .QN());
   DFF_X1 \buffer_reg[0][2][2][10]  (.D(\input_filter[2][2] [10]), .CK(n_55_12), 
      .Q(\buffer[0][2][2] [10]), .QN());
   DFF_X1 \buffer_reg[0][2][2][9]  (.D(\input_filter[2][2] [9]), .CK(n_55_12), 
      .Q(\buffer[0][2][2] [9]), .QN());
   DFF_X1 \buffer_reg[0][2][2][8]  (.D(\input_filter[2][2] [8]), .CK(n_55_12), 
      .Q(\buffer[0][2][2] [8]), .QN());
   DFF_X1 \buffer_reg[0][2][2][7]  (.D(\input_filter[2][2] [7]), .CK(n_55_12), 
      .Q(\buffer[0][2][2] [7]), .QN());
   DFF_X1 \buffer_reg[0][2][2][6]  (.D(\input_filter[2][2] [6]), .CK(n_55_12), 
      .Q(\buffer[0][2][2] [6]), .QN());
   DFF_X1 \buffer_reg[0][2][2][5]  (.D(\input_filter[2][2] [5]), .CK(n_55_12), 
      .Q(\buffer[0][2][2] [5]), .QN());
   DFF_X1 \buffer_reg[0][2][2][4]  (.D(\input_filter[2][2] [4]), .CK(n_55_12), 
      .Q(\buffer[0][2][2] [4]), .QN());
   DFF_X1 \buffer_reg[0][2][2][3]  (.D(\input_filter[2][2] [3]), .CK(n_55_12), 
      .Q(\buffer[0][2][2] [3]), .QN());
   DFF_X1 \buffer_reg[0][2][2][2]  (.D(\input_filter[2][2] [2]), .CK(n_55_12), 
      .Q(\buffer[0][2][2] [2]), .QN());
   DFF_X1 \buffer_reg[0][2][2][1]  (.D(\input_filter[2][2] [1]), .CK(n_55_12), 
      .Q(\buffer[0][2][2] [1]), .QN());
   DFF_X1 \buffer_reg[0][2][2][0]  (.D(\input_filter[2][2] [0]), .CK(n_55_12), 
      .Q(\buffer[0][2][2] [0]), .QN());
   DFF_X1 \buffer_reg[0][0][0][15]  (.D(\input_filter[0][0] [15]), .CK(n_55_12), 
      .Q(\buffer[0][0][0] [15]), .QN());
   DFF_X1 \buffer_reg[0][0][0][14]  (.D(\input_filter[0][0] [14]), .CK(n_55_12), 
      .Q(\buffer[0][0][0] [14]), .QN());
   DFF_X1 \buffer_reg[0][0][0][13]  (.D(\input_filter[0][0] [13]), .CK(n_55_12), 
      .Q(\buffer[0][0][0] [13]), .QN());
   DFF_X1 \buffer_reg[0][0][0][12]  (.D(\input_filter[0][0] [12]), .CK(n_55_12), 
      .Q(\buffer[0][0][0] [12]), .QN());
   DFF_X1 \buffer_reg[0][0][0][11]  (.D(\input_filter[0][0] [11]), .CK(n_55_12), 
      .Q(\buffer[0][0][0] [11]), .QN());
   DFF_X1 \buffer_reg[0][0][0][10]  (.D(\input_filter[0][0] [10]), .CK(n_55_12), 
      .Q(\buffer[0][0][0] [10]), .QN());
   DFF_X1 \buffer_reg[0][0][0][9]  (.D(\input_filter[0][0] [9]), .CK(n_55_12), 
      .Q(\buffer[0][0][0] [9]), .QN());
   DFF_X1 \buffer_reg[0][0][0][8]  (.D(\input_filter[0][0] [8]), .CK(n_55_12), 
      .Q(\buffer[0][0][0] [8]), .QN());
   DFF_X1 \buffer_reg[0][0][0][7]  (.D(\input_filter[0][0] [7]), .CK(n_55_12), 
      .Q(\buffer[0][0][0] [7]), .QN());
   DFF_X1 \buffer_reg[0][0][0][6]  (.D(\input_filter[0][0] [6]), .CK(n_55_12), 
      .Q(\buffer[0][0][0] [6]), .QN());
   DFF_X1 \buffer_reg[0][0][0][5]  (.D(\input_filter[0][0] [5]), .CK(n_55_12), 
      .Q(\buffer[0][0][0] [5]), .QN());
   DFF_X1 \buffer_reg[0][0][0][4]  (.D(\input_filter[0][0] [4]), .CK(n_55_12), 
      .Q(\buffer[0][0][0] [4]), .QN());
   DFF_X1 \buffer_reg[0][0][0][3]  (.D(\input_filter[0][0] [3]), .CK(n_55_12), 
      .Q(\buffer[0][0][0] [3]), .QN());
   DFF_X1 \buffer_reg[0][0][0][2]  (.D(\input_filter[0][0] [2]), .CK(n_55_12), 
      .Q(\buffer[0][0][0] [2]), .QN());
   DFF_X1 \buffer_reg[0][0][0][1]  (.D(\input_filter[0][0] [1]), .CK(n_55_12), 
      .Q(\buffer[0][0][0] [1]), .QN());
   DFF_X1 \buffer_reg[0][0][0][0]  (.D(\input_filter[0][0] [0]), .CK(n_55_12), 
      .Q(\buffer[0][0][0] [0]), .QN());
   DFF_X1 \buffer_reg[13][3][2][15]  (.D(\input_filter[3][2] [15]), .CK(n_55_15), 
      .Q(\buffer[13][3][2] [15]), .QN());
   DFF_X1 \buffer_reg[13][3][2][14]  (.D(\input_filter[3][2] [14]), .CK(n_55_15), 
      .Q(\buffer[13][3][2] [14]), .QN());
   DFF_X1 \buffer_reg[13][3][2][13]  (.D(\input_filter[3][2] [13]), .CK(n_55_15), 
      .Q(\buffer[13][3][2] [13]), .QN());
   DFF_X1 \buffer_reg[13][3][2][12]  (.D(\input_filter[3][2] [12]), .CK(n_55_15), 
      .Q(\buffer[13][3][2] [12]), .QN());
   DFF_X1 \buffer_reg[13][3][2][11]  (.D(\input_filter[3][2] [11]), .CK(n_55_15), 
      .Q(\buffer[13][3][2] [11]), .QN());
   DFF_X1 \buffer_reg[13][3][2][10]  (.D(\input_filter[3][2] [10]), .CK(n_55_15), 
      .Q(\buffer[13][3][2] [10]), .QN());
   DFF_X1 \buffer_reg[13][3][2][9]  (.D(\input_filter[3][2] [9]), .CK(n_55_15), 
      .Q(\buffer[13][3][2] [9]), .QN());
   DFF_X1 \buffer_reg[13][3][2][8]  (.D(\input_filter[3][2] [8]), .CK(n_55_15), 
      .Q(\buffer[13][3][2] [8]), .QN());
   DFF_X1 \buffer_reg[13][3][2][7]  (.D(\input_filter[3][2] [7]), .CK(n_55_15), 
      .Q(\buffer[13][3][2] [7]), .QN());
   DFF_X1 \buffer_reg[13][3][2][6]  (.D(\input_filter[3][2] [6]), .CK(n_55_15), 
      .Q(\buffer[13][3][2] [6]), .QN());
   DFF_X1 \buffer_reg[13][3][2][5]  (.D(\input_filter[3][2] [5]), .CK(n_55_15), 
      .Q(\buffer[13][3][2] [5]), .QN());
   DFF_X1 \buffer_reg[13][3][2][4]  (.D(\input_filter[3][2] [4]), .CK(n_55_15), 
      .Q(\buffer[13][3][2] [4]), .QN());
   DFF_X1 \buffer_reg[13][3][2][3]  (.D(\input_filter[3][2] [3]), .CK(n_55_15), 
      .Q(\buffer[13][3][2] [3]), .QN());
   DFF_X1 \buffer_reg[13][3][2][2]  (.D(\input_filter[3][2] [2]), .CK(n_55_15), 
      .Q(\buffer[13][3][2] [2]), .QN());
   DFF_X1 \buffer_reg[13][3][2][1]  (.D(\input_filter[3][2] [1]), .CK(n_55_15), 
      .Q(\buffer[13][3][2] [1]), .QN());
   DFF_X1 \buffer_reg[13][3][2][0]  (.D(\input_filter[3][2] [0]), .CK(n_55_15), 
      .Q(\buffer[13][3][2] [0]), .QN());
   DFF_X1 \buffer_reg[14][3][2][15]  (.D(\input_filter[3][2] [15]), .CK(n_55_14), 
      .Q(\buffer[14][3][2] [15]), .QN());
   DFF_X1 \buffer_reg[14][3][2][14]  (.D(\input_filter[3][2] [14]), .CK(n_55_14), 
      .Q(\buffer[14][3][2] [14]), .QN());
   DFF_X1 \buffer_reg[14][3][2][13]  (.D(\input_filter[3][2] [13]), .CK(n_55_14), 
      .Q(\buffer[14][3][2] [13]), .QN());
   DFF_X1 \buffer_reg[14][3][2][12]  (.D(\input_filter[3][2] [12]), .CK(n_55_14), 
      .Q(\buffer[14][3][2] [12]), .QN());
   DFF_X1 \buffer_reg[14][3][2][11]  (.D(\input_filter[3][2] [11]), .CK(n_55_14), 
      .Q(\buffer[14][3][2] [11]), .QN());
   DFF_X1 \buffer_reg[14][3][2][10]  (.D(\input_filter[3][2] [10]), .CK(n_55_14), 
      .Q(\buffer[14][3][2] [10]), .QN());
   DFF_X1 \buffer_reg[14][3][2][9]  (.D(\input_filter[3][2] [9]), .CK(n_55_14), 
      .Q(\buffer[14][3][2] [9]), .QN());
   DFF_X1 \buffer_reg[14][3][2][8]  (.D(\input_filter[3][2] [8]), .CK(n_55_14), 
      .Q(\buffer[14][3][2] [8]), .QN());
   DFF_X1 \buffer_reg[14][3][2][7]  (.D(\input_filter[3][2] [7]), .CK(n_55_14), 
      .Q(\buffer[14][3][2] [7]), .QN());
   DFF_X1 \buffer_reg[14][3][2][6]  (.D(\input_filter[3][2] [6]), .CK(n_55_14), 
      .Q(\buffer[14][3][2] [6]), .QN());
   DFF_X1 \buffer_reg[14][3][2][5]  (.D(\input_filter[3][2] [5]), .CK(n_55_14), 
      .Q(\buffer[14][3][2] [5]), .QN());
   DFF_X1 \buffer_reg[14][3][2][4]  (.D(\input_filter[3][2] [4]), .CK(n_55_14), 
      .Q(\buffer[14][3][2] [4]), .QN());
   DFF_X1 \buffer_reg[14][3][2][3]  (.D(\input_filter[3][2] [3]), .CK(n_55_14), 
      .Q(\buffer[14][3][2] [3]), .QN());
   DFF_X1 \buffer_reg[14][3][2][2]  (.D(\input_filter[3][2] [2]), .CK(n_55_14), 
      .Q(\buffer[14][3][2] [2]), .QN());
   DFF_X1 \buffer_reg[14][3][2][1]  (.D(\input_filter[3][2] [1]), .CK(n_55_14), 
      .Q(\buffer[14][3][2] [1]), .QN());
   DFF_X1 \buffer_reg[14][3][2][0]  (.D(\input_filter[3][2] [0]), .CK(n_55_14), 
      .Q(\buffer[14][3][2] [0]), .QN());
   DFF_X1 \buffer_reg[15][3][2][15]  (.D(\input_filter[3][2] [15]), .CK(n_55_13), 
      .Q(\buffer[15][3][2] [15]), .QN());
   DFF_X1 \buffer_reg[15][3][2][14]  (.D(\input_filter[3][2] [14]), .CK(n_55_13), 
      .Q(\buffer[15][3][2] [14]), .QN());
   DFF_X1 \buffer_reg[15][3][2][13]  (.D(\input_filter[3][2] [13]), .CK(n_55_13), 
      .Q(\buffer[15][3][2] [13]), .QN());
   DFF_X1 \buffer_reg[15][3][2][12]  (.D(\input_filter[3][2] [12]), .CK(n_55_13), 
      .Q(\buffer[15][3][2] [12]), .QN());
   DFF_X1 \buffer_reg[15][3][2][11]  (.D(\input_filter[3][2] [11]), .CK(n_55_13), 
      .Q(\buffer[15][3][2] [11]), .QN());
   DFF_X1 \buffer_reg[15][3][2][10]  (.D(\input_filter[3][2] [10]), .CK(n_55_13), 
      .Q(\buffer[15][3][2] [10]), .QN());
   DFF_X1 \buffer_reg[15][3][2][9]  (.D(\input_filter[3][2] [9]), .CK(n_55_13), 
      .Q(\buffer[15][3][2] [9]), .QN());
   DFF_X1 \buffer_reg[15][3][2][8]  (.D(\input_filter[3][2] [8]), .CK(n_55_13), 
      .Q(\buffer[15][3][2] [8]), .QN());
   DFF_X1 \buffer_reg[15][3][2][7]  (.D(\input_filter[3][2] [7]), .CK(n_55_13), 
      .Q(\buffer[15][3][2] [7]), .QN());
   DFF_X1 \buffer_reg[15][3][2][6]  (.D(\input_filter[3][2] [6]), .CK(n_55_13), 
      .Q(\buffer[15][3][2] [6]), .QN());
   DFF_X1 \buffer_reg[15][3][2][5]  (.D(\input_filter[3][2] [5]), .CK(n_55_13), 
      .Q(\buffer[15][3][2] [5]), .QN());
   DFF_X1 \buffer_reg[15][3][2][4]  (.D(\input_filter[3][2] [4]), .CK(n_55_13), 
      .Q(\buffer[15][3][2] [4]), .QN());
   DFF_X1 \buffer_reg[15][3][2][3]  (.D(\input_filter[3][2] [3]), .CK(n_55_13), 
      .Q(\buffer[15][3][2] [3]), .QN());
   DFF_X1 \buffer_reg[15][3][2][2]  (.D(\input_filter[3][2] [2]), .CK(n_55_13), 
      .Q(\buffer[15][3][2] [2]), .QN());
   DFF_X1 \buffer_reg[15][3][2][1]  (.D(\input_filter[3][2] [1]), .CK(n_55_13), 
      .Q(\buffer[15][3][2] [1]), .QN());
   DFF_X1 \buffer_reg[15][3][2][0]  (.D(\input_filter[3][2] [0]), .CK(n_55_13), 
      .Q(\buffer[15][3][2] [0]), .QN());
   CLKGATETST_X1 \clk_gate_buffer_reg[12][3][2]_reg  (.CK(read), .E(n_12), 
      .SE(1'b0), .GCK(n_55_0));
   CLKGATETST_X1 \clk_gate_buffer_reg[11][3][2]_reg  (.CK(read), .E(n_11), 
      .SE(1'b0), .GCK(n_55_1));
   CLKGATETST_X1 \clk_gate_buffer_reg[10][3][2]_reg  (.CK(read), .E(n_10), 
      .SE(1'b0), .GCK(n_55_2));
   CLKGATETST_X1 \clk_gate_buffer_reg[9][3][2]_reg  (.CK(read), .E(n_9), 
      .SE(1'b0), .GCK(n_55_3));
   CLKGATETST_X1 \clk_gate_buffer_reg[8][3][2]_reg  (.CK(read), .E(n_8), 
      .SE(1'b0), .GCK(n_55_4));
   CLKGATETST_X1 \clk_gate_buffer_reg[7][3][2]_reg  (.CK(read), .E(n_7), 
      .SE(1'b0), .GCK(n_55_5));
   CLKGATETST_X1 \clk_gate_buffer_reg[6][3][2]_reg  (.CK(read), .E(n_6), 
      .SE(1'b0), .GCK(n_55_6));
   CLKGATETST_X1 \clk_gate_buffer_reg[5][3][2]_reg  (.CK(read), .E(n_5), 
      .SE(1'b0), .GCK(n_55_7));
   CLKGATETST_X1 \clk_gate_buffer_reg[4][3][2]_reg  (.CK(read), .E(n_4), 
      .SE(1'b0), .GCK(n_55_8));
   CLKGATETST_X1 \clk_gate_buffer_reg[3][3][2]_reg  (.CK(read), .E(n_3), 
      .SE(1'b0), .GCK(n_55_9));
   CLKGATETST_X1 \clk_gate_buffer_reg[2][3][2]_reg  (.CK(read), .E(n_2), 
      .SE(1'b0), .GCK(n_55_10));
   CLKGATETST_X1 \clk_gate_buffer_reg[1][3][2]_reg  (.CK(read), .E(n_1), 
      .SE(1'b0), .GCK(n_55_11));
   CLKGATETST_X1 \clk_gate_buffer_reg[0][3][2]_reg  (.CK(read), .E(n_0), 
      .SE(1'b0), .GCK(n_55_12));
   CLKGATETST_X1 \clk_gate_buffer_reg[15][3][1]_reg  (.CK(read), .E(n_15), 
      .SE(1'b0), .GCK(n_55_13));
   CLKGATETST_X1 \clk_gate_buffer_reg[14][3][1]_reg  (.CK(read), .E(n_14), 
      .SE(1'b0), .GCK(n_55_14));
   CLKGATETST_X1 \clk_gate_buffer_reg[13][3][1]_reg  (.CK(read), .E(n_13), 
      .SE(1'b0), .GCK(n_55_15));
   DFF_X1 \buffer_reg[3][0][0][15]  (.D(\input_filter[0][0] [15]), .CK(n_56_0), 
      .Q(\buffer[3][0][0] [15]), .QN());
   DFF_X1 \buffer_reg[3][0][0][14]  (.D(\input_filter[0][0] [14]), .CK(n_56_0), 
      .Q(\buffer[3][0][0] [14]), .QN());
   DFF_X1 \buffer_reg[3][0][0][13]  (.D(\input_filter[0][0] [13]), .CK(n_56_0), 
      .Q(\buffer[3][0][0] [13]), .QN());
   DFF_X1 \buffer_reg[3][0][0][12]  (.D(\input_filter[0][0] [12]), .CK(n_56_0), 
      .Q(\buffer[3][0][0] [12]), .QN());
   DFF_X1 \buffer_reg[3][0][0][11]  (.D(\input_filter[0][0] [11]), .CK(n_56_0), 
      .Q(\buffer[3][0][0] [11]), .QN());
   DFF_X1 \buffer_reg[3][0][0][10]  (.D(\input_filter[0][0] [10]), .CK(n_56_0), 
      .Q(\buffer[3][0][0] [10]), .QN());
   DFF_X1 \buffer_reg[3][0][0][9]  (.D(\input_filter[0][0] [9]), .CK(n_56_0), 
      .Q(\buffer[3][0][0] [9]), .QN());
   DFF_X1 \buffer_reg[3][0][0][8]  (.D(\input_filter[0][0] [8]), .CK(n_56_0), 
      .Q(\buffer[3][0][0] [8]), .QN());
   DFF_X1 \buffer_reg[3][0][0][7]  (.D(\input_filter[0][0] [7]), .CK(n_56_0), 
      .Q(\buffer[3][0][0] [7]), .QN());
   DFF_X1 \buffer_reg[3][0][0][6]  (.D(\input_filter[0][0] [6]), .CK(n_56_0), 
      .Q(\buffer[3][0][0] [6]), .QN());
   DFF_X1 \buffer_reg[3][0][0][5]  (.D(\input_filter[0][0] [5]), .CK(n_56_0), 
      .Q(\buffer[3][0][0] [5]), .QN());
   DFF_X1 \buffer_reg[3][0][0][4]  (.D(\input_filter[0][0] [4]), .CK(n_56_0), 
      .Q(\buffer[3][0][0] [4]), .QN());
   DFF_X1 \buffer_reg[3][0][0][3]  (.D(\input_filter[0][0] [3]), .CK(n_56_0), 
      .Q(\buffer[3][0][0] [3]), .QN());
   DFF_X1 \buffer_reg[3][0][0][2]  (.D(\input_filter[0][0] [2]), .CK(n_56_0), 
      .Q(\buffer[3][0][0] [2]), .QN());
   DFF_X1 \buffer_reg[3][0][0][1]  (.D(\input_filter[0][0] [1]), .CK(n_56_0), 
      .Q(\buffer[3][0][0] [1]), .QN());
   DFF_X1 \buffer_reg[3][0][0][0]  (.D(\input_filter[0][0] [0]), .CK(n_56_0), 
      .Q(\buffer[3][0][0] [0]), .QN());
   DFF_X1 \buffer_reg[4][0][0][15]  (.D(\input_filter[0][0] [15]), .CK(n_56_1), 
      .Q(\buffer[4][0][0] [15]), .QN());
   DFF_X1 \buffer_reg[4][0][0][14]  (.D(\input_filter[0][0] [14]), .CK(n_56_1), 
      .Q(\buffer[4][0][0] [14]), .QN());
   DFF_X1 \buffer_reg[4][0][0][13]  (.D(\input_filter[0][0] [13]), .CK(n_56_1), 
      .Q(\buffer[4][0][0] [13]), .QN());
   DFF_X1 \buffer_reg[4][0][0][12]  (.D(\input_filter[0][0] [12]), .CK(n_56_1), 
      .Q(\buffer[4][0][0] [12]), .QN());
   DFF_X1 \buffer_reg[4][0][0][11]  (.D(\input_filter[0][0] [11]), .CK(n_56_1), 
      .Q(\buffer[4][0][0] [11]), .QN());
   DFF_X1 \buffer_reg[4][0][0][10]  (.D(\input_filter[0][0] [10]), .CK(n_56_1), 
      .Q(\buffer[4][0][0] [10]), .QN());
   DFF_X1 \buffer_reg[4][0][0][9]  (.D(\input_filter[0][0] [9]), .CK(n_56_1), 
      .Q(\buffer[4][0][0] [9]), .QN());
   DFF_X1 \buffer_reg[4][0][0][8]  (.D(\input_filter[0][0] [8]), .CK(n_56_1), 
      .Q(\buffer[4][0][0] [8]), .QN());
   DFF_X1 \buffer_reg[4][0][0][7]  (.D(\input_filter[0][0] [7]), .CK(n_56_1), 
      .Q(\buffer[4][0][0] [7]), .QN());
   DFF_X1 \buffer_reg[4][0][0][6]  (.D(\input_filter[0][0] [6]), .CK(n_56_1), 
      .Q(\buffer[4][0][0] [6]), .QN());
   DFF_X1 \buffer_reg[4][0][0][5]  (.D(\input_filter[0][0] [5]), .CK(n_56_1), 
      .Q(\buffer[4][0][0] [5]), .QN());
   DFF_X1 \buffer_reg[4][0][0][4]  (.D(\input_filter[0][0] [4]), .CK(n_56_1), 
      .Q(\buffer[4][0][0] [4]), .QN());
   DFF_X1 \buffer_reg[4][0][0][3]  (.D(\input_filter[0][0] [3]), .CK(n_56_1), 
      .Q(\buffer[4][0][0] [3]), .QN());
   DFF_X1 \buffer_reg[4][0][0][2]  (.D(\input_filter[0][0] [2]), .CK(n_56_1), 
      .Q(\buffer[4][0][0] [2]), .QN());
   DFF_X1 \buffer_reg[4][0][0][1]  (.D(\input_filter[0][0] [1]), .CK(n_56_1), 
      .Q(\buffer[4][0][0] [1]), .QN());
   DFF_X1 \buffer_reg[4][0][0][0]  (.D(\input_filter[0][0] [0]), .CK(n_56_1), 
      .Q(\buffer[4][0][0] [0]), .QN());
   DFF_X1 \buffer_reg[5][0][0][15]  (.D(\input_filter[0][0] [15]), .CK(n_56_2), 
      .Q(\buffer[5][0][0] [15]), .QN());
   DFF_X1 \buffer_reg[5][0][0][14]  (.D(\input_filter[0][0] [14]), .CK(n_56_2), 
      .Q(\buffer[5][0][0] [14]), .QN());
   DFF_X1 \buffer_reg[5][0][0][13]  (.D(\input_filter[0][0] [13]), .CK(n_56_2), 
      .Q(\buffer[5][0][0] [13]), .QN());
   DFF_X1 \buffer_reg[5][0][0][12]  (.D(\input_filter[0][0] [12]), .CK(n_56_2), 
      .Q(\buffer[5][0][0] [12]), .QN());
   DFF_X1 \buffer_reg[5][0][0][11]  (.D(\input_filter[0][0] [11]), .CK(n_56_2), 
      .Q(\buffer[5][0][0] [11]), .QN());
   DFF_X1 \buffer_reg[5][0][0][10]  (.D(\input_filter[0][0] [10]), .CK(n_56_2), 
      .Q(\buffer[5][0][0] [10]), .QN());
   DFF_X1 \buffer_reg[5][0][0][9]  (.D(\input_filter[0][0] [9]), .CK(n_56_2), 
      .Q(\buffer[5][0][0] [9]), .QN());
   DFF_X1 \buffer_reg[5][0][0][8]  (.D(\input_filter[0][0] [8]), .CK(n_56_2), 
      .Q(\buffer[5][0][0] [8]), .QN());
   DFF_X1 \buffer_reg[5][0][0][7]  (.D(\input_filter[0][0] [7]), .CK(n_56_2), 
      .Q(\buffer[5][0][0] [7]), .QN());
   DFF_X1 \buffer_reg[5][0][0][6]  (.D(\input_filter[0][0] [6]), .CK(n_56_2), 
      .Q(\buffer[5][0][0] [6]), .QN());
   DFF_X1 \buffer_reg[5][0][0][5]  (.D(\input_filter[0][0] [5]), .CK(n_56_2), 
      .Q(\buffer[5][0][0] [5]), .QN());
   DFF_X1 \buffer_reg[5][0][0][4]  (.D(\input_filter[0][0] [4]), .CK(n_56_2), 
      .Q(\buffer[5][0][0] [4]), .QN());
   DFF_X1 \buffer_reg[5][0][0][3]  (.D(\input_filter[0][0] [3]), .CK(n_56_2), 
      .Q(\buffer[5][0][0] [3]), .QN());
   DFF_X1 \buffer_reg[5][0][0][2]  (.D(\input_filter[0][0] [2]), .CK(n_56_2), 
      .Q(\buffer[5][0][0] [2]), .QN());
   DFF_X1 \buffer_reg[5][0][0][1]  (.D(\input_filter[0][0] [1]), .CK(n_56_2), 
      .Q(\buffer[5][0][0] [1]), .QN());
   DFF_X1 \buffer_reg[5][0][0][0]  (.D(\input_filter[0][0] [0]), .CK(n_56_2), 
      .Q(\buffer[5][0][0] [0]), .QN());
   DFF_X1 \buffer_reg[6][0][0][15]  (.D(\input_filter[0][0] [15]), .CK(n_56_3), 
      .Q(\buffer[6][0][0] [15]), .QN());
   DFF_X1 \buffer_reg[6][0][0][14]  (.D(\input_filter[0][0] [14]), .CK(n_56_3), 
      .Q(\buffer[6][0][0] [14]), .QN());
   DFF_X1 \buffer_reg[6][0][0][13]  (.D(\input_filter[0][0] [13]), .CK(n_56_3), 
      .Q(\buffer[6][0][0] [13]), .QN());
   DFF_X1 \buffer_reg[6][0][0][12]  (.D(\input_filter[0][0] [12]), .CK(n_56_3), 
      .Q(\buffer[6][0][0] [12]), .QN());
   DFF_X1 \buffer_reg[6][0][0][11]  (.D(\input_filter[0][0] [11]), .CK(n_56_3), 
      .Q(\buffer[6][0][0] [11]), .QN());
   DFF_X1 \buffer_reg[6][0][0][10]  (.D(\input_filter[0][0] [10]), .CK(n_56_3), 
      .Q(\buffer[6][0][0] [10]), .QN());
   DFF_X1 \buffer_reg[6][0][0][9]  (.D(\input_filter[0][0] [9]), .CK(n_56_3), 
      .Q(\buffer[6][0][0] [9]), .QN());
   DFF_X1 \buffer_reg[6][0][0][8]  (.D(\input_filter[0][0] [8]), .CK(n_56_3), 
      .Q(\buffer[6][0][0] [8]), .QN());
   DFF_X1 \buffer_reg[6][0][0][7]  (.D(\input_filter[0][0] [7]), .CK(n_56_3), 
      .Q(\buffer[6][0][0] [7]), .QN());
   DFF_X1 \buffer_reg[6][0][0][6]  (.D(\input_filter[0][0] [6]), .CK(n_56_3), 
      .Q(\buffer[6][0][0] [6]), .QN());
   DFF_X1 \buffer_reg[6][0][0][5]  (.D(\input_filter[0][0] [5]), .CK(n_56_3), 
      .Q(\buffer[6][0][0] [5]), .QN());
   DFF_X1 \buffer_reg[6][0][0][4]  (.D(\input_filter[0][0] [4]), .CK(n_56_3), 
      .Q(\buffer[6][0][0] [4]), .QN());
   DFF_X1 \buffer_reg[6][0][0][3]  (.D(\input_filter[0][0] [3]), .CK(n_56_3), 
      .Q(\buffer[6][0][0] [3]), .QN());
   DFF_X1 \buffer_reg[6][0][0][2]  (.D(\input_filter[0][0] [2]), .CK(n_56_3), 
      .Q(\buffer[6][0][0] [2]), .QN());
   DFF_X1 \buffer_reg[6][0][0][1]  (.D(\input_filter[0][0] [1]), .CK(n_56_3), 
      .Q(\buffer[6][0][0] [1]), .QN());
   DFF_X1 \buffer_reg[6][0][0][0]  (.D(\input_filter[0][0] [0]), .CK(n_56_3), 
      .Q(\buffer[6][0][0] [0]), .QN());
   DFF_X1 \buffer_reg[7][0][0][15]  (.D(\input_filter[0][0] [15]), .CK(n_56_4), 
      .Q(\buffer[7][0][0] [15]), .QN());
   DFF_X1 \buffer_reg[7][0][0][14]  (.D(\input_filter[0][0] [14]), .CK(n_56_4), 
      .Q(\buffer[7][0][0] [14]), .QN());
   DFF_X1 \buffer_reg[7][0][0][13]  (.D(\input_filter[0][0] [13]), .CK(n_56_4), 
      .Q(\buffer[7][0][0] [13]), .QN());
   DFF_X1 \buffer_reg[7][0][0][12]  (.D(\input_filter[0][0] [12]), .CK(n_56_4), 
      .Q(\buffer[7][0][0] [12]), .QN());
   DFF_X1 \buffer_reg[7][0][0][11]  (.D(\input_filter[0][0] [11]), .CK(n_56_4), 
      .Q(\buffer[7][0][0] [11]), .QN());
   DFF_X1 \buffer_reg[7][0][0][10]  (.D(\input_filter[0][0] [10]), .CK(n_56_4), 
      .Q(\buffer[7][0][0] [10]), .QN());
   DFF_X1 \buffer_reg[7][0][0][9]  (.D(\input_filter[0][0] [9]), .CK(n_56_4), 
      .Q(\buffer[7][0][0] [9]), .QN());
   DFF_X1 \buffer_reg[7][0][0][8]  (.D(\input_filter[0][0] [8]), .CK(n_56_4), 
      .Q(\buffer[7][0][0] [8]), .QN());
   DFF_X1 \buffer_reg[7][0][0][7]  (.D(\input_filter[0][0] [7]), .CK(n_56_4), 
      .Q(\buffer[7][0][0] [7]), .QN());
   DFF_X1 \buffer_reg[7][0][0][6]  (.D(\input_filter[0][0] [6]), .CK(n_56_4), 
      .Q(\buffer[7][0][0] [6]), .QN());
   DFF_X1 \buffer_reg[7][0][0][5]  (.D(\input_filter[0][0] [5]), .CK(n_56_4), 
      .Q(\buffer[7][0][0] [5]), .QN());
   DFF_X1 \buffer_reg[7][0][0][4]  (.D(\input_filter[0][0] [4]), .CK(n_56_4), 
      .Q(\buffer[7][0][0] [4]), .QN());
   DFF_X1 \buffer_reg[7][0][0][3]  (.D(\input_filter[0][0] [3]), .CK(n_56_4), 
      .Q(\buffer[7][0][0] [3]), .QN());
   DFF_X1 \buffer_reg[7][0][0][2]  (.D(\input_filter[0][0] [2]), .CK(n_56_4), 
      .Q(\buffer[7][0][0] [2]), .QN());
   DFF_X1 \buffer_reg[7][0][0][1]  (.D(\input_filter[0][0] [1]), .CK(n_56_4), 
      .Q(\buffer[7][0][0] [1]), .QN());
   DFF_X1 \buffer_reg[7][0][0][0]  (.D(\input_filter[0][0] [0]), .CK(n_56_4), 
      .Q(\buffer[7][0][0] [0]), .QN());
   DFF_X1 \buffer_reg[8][0][0][15]  (.D(\input_filter[0][0] [15]), .CK(n_56_5), 
      .Q(\buffer[8][0][0] [15]), .QN());
   DFF_X1 \buffer_reg[8][0][0][14]  (.D(\input_filter[0][0] [14]), .CK(n_56_5), 
      .Q(\buffer[8][0][0] [14]), .QN());
   DFF_X1 \buffer_reg[8][0][0][13]  (.D(\input_filter[0][0] [13]), .CK(n_56_5), 
      .Q(\buffer[8][0][0] [13]), .QN());
   DFF_X1 \buffer_reg[8][0][0][12]  (.D(\input_filter[0][0] [12]), .CK(n_56_5), 
      .Q(\buffer[8][0][0] [12]), .QN());
   DFF_X1 \buffer_reg[8][0][0][11]  (.D(\input_filter[0][0] [11]), .CK(n_56_5), 
      .Q(\buffer[8][0][0] [11]), .QN());
   DFF_X1 \buffer_reg[8][0][0][10]  (.D(\input_filter[0][0] [10]), .CK(n_56_5), 
      .Q(\buffer[8][0][0] [10]), .QN());
   DFF_X1 \buffer_reg[8][0][0][9]  (.D(\input_filter[0][0] [9]), .CK(n_56_5), 
      .Q(\buffer[8][0][0] [9]), .QN());
   DFF_X1 \buffer_reg[8][0][0][8]  (.D(\input_filter[0][0] [8]), .CK(n_56_5), 
      .Q(\buffer[8][0][0] [8]), .QN());
   DFF_X1 \buffer_reg[8][0][0][7]  (.D(\input_filter[0][0] [7]), .CK(n_56_5), 
      .Q(\buffer[8][0][0] [7]), .QN());
   DFF_X1 \buffer_reg[8][0][0][6]  (.D(\input_filter[0][0] [6]), .CK(n_56_5), 
      .Q(\buffer[8][0][0] [6]), .QN());
   DFF_X1 \buffer_reg[8][0][0][5]  (.D(\input_filter[0][0] [5]), .CK(n_56_5), 
      .Q(\buffer[8][0][0] [5]), .QN());
   DFF_X1 \buffer_reg[8][0][0][4]  (.D(\input_filter[0][0] [4]), .CK(n_56_5), 
      .Q(\buffer[8][0][0] [4]), .QN());
   DFF_X1 \buffer_reg[8][0][0][3]  (.D(\input_filter[0][0] [3]), .CK(n_56_5), 
      .Q(\buffer[8][0][0] [3]), .QN());
   DFF_X1 \buffer_reg[8][0][0][2]  (.D(\input_filter[0][0] [2]), .CK(n_56_5), 
      .Q(\buffer[8][0][0] [2]), .QN());
   DFF_X1 \buffer_reg[8][0][0][1]  (.D(\input_filter[0][0] [1]), .CK(n_56_5), 
      .Q(\buffer[8][0][0] [1]), .QN());
   DFF_X1 \buffer_reg[8][0][0][0]  (.D(\input_filter[0][0] [0]), .CK(n_56_5), 
      .Q(\buffer[8][0][0] [0]), .QN());
   DFF_X1 \buffer_reg[9][0][0][15]  (.D(\input_filter[0][0] [15]), .CK(n_56_6), 
      .Q(\buffer[9][0][0] [15]), .QN());
   DFF_X1 \buffer_reg[9][0][0][14]  (.D(\input_filter[0][0] [14]), .CK(n_56_6), 
      .Q(\buffer[9][0][0] [14]), .QN());
   DFF_X1 \buffer_reg[9][0][0][13]  (.D(\input_filter[0][0] [13]), .CK(n_56_6), 
      .Q(\buffer[9][0][0] [13]), .QN());
   DFF_X1 \buffer_reg[9][0][0][12]  (.D(\input_filter[0][0] [12]), .CK(n_56_6), 
      .Q(\buffer[9][0][0] [12]), .QN());
   DFF_X1 \buffer_reg[9][0][0][11]  (.D(\input_filter[0][0] [11]), .CK(n_56_6), 
      .Q(\buffer[9][0][0] [11]), .QN());
   DFF_X1 \buffer_reg[9][0][0][10]  (.D(\input_filter[0][0] [10]), .CK(n_56_6), 
      .Q(\buffer[9][0][0] [10]), .QN());
   DFF_X1 \buffer_reg[9][0][0][9]  (.D(\input_filter[0][0] [9]), .CK(n_56_6), 
      .Q(\buffer[9][0][0] [9]), .QN());
   DFF_X1 \buffer_reg[9][0][0][8]  (.D(\input_filter[0][0] [8]), .CK(n_56_6), 
      .Q(\buffer[9][0][0] [8]), .QN());
   DFF_X1 \buffer_reg[9][0][0][7]  (.D(\input_filter[0][0] [7]), .CK(n_56_6), 
      .Q(\buffer[9][0][0] [7]), .QN());
   DFF_X1 \buffer_reg[9][0][0][6]  (.D(\input_filter[0][0] [6]), .CK(n_56_6), 
      .Q(\buffer[9][0][0] [6]), .QN());
   DFF_X1 \buffer_reg[9][0][0][5]  (.D(\input_filter[0][0] [5]), .CK(n_56_6), 
      .Q(\buffer[9][0][0] [5]), .QN());
   DFF_X1 \buffer_reg[9][0][0][4]  (.D(\input_filter[0][0] [4]), .CK(n_56_6), 
      .Q(\buffer[9][0][0] [4]), .QN());
   DFF_X1 \buffer_reg[9][0][0][3]  (.D(\input_filter[0][0] [3]), .CK(n_56_6), 
      .Q(\buffer[9][0][0] [3]), .QN());
   DFF_X1 \buffer_reg[9][0][0][2]  (.D(\input_filter[0][0] [2]), .CK(n_56_6), 
      .Q(\buffer[9][0][0] [2]), .QN());
   DFF_X1 \buffer_reg[9][0][0][1]  (.D(\input_filter[0][0] [1]), .CK(n_56_6), 
      .Q(\buffer[9][0][0] [1]), .QN());
   DFF_X1 \buffer_reg[9][0][0][0]  (.D(\input_filter[0][0] [0]), .CK(n_56_6), 
      .Q(\buffer[9][0][0] [0]), .QN());
   DFF_X1 \buffer_reg[10][0][0][15]  (.D(\input_filter[0][0] [15]), .CK(n_56_7), 
      .Q(\buffer[10][0][0] [15]), .QN());
   DFF_X1 \buffer_reg[10][0][0][14]  (.D(\input_filter[0][0] [14]), .CK(n_56_7), 
      .Q(\buffer[10][0][0] [14]), .QN());
   DFF_X1 \buffer_reg[10][0][0][13]  (.D(\input_filter[0][0] [13]), .CK(n_56_7), 
      .Q(\buffer[10][0][0] [13]), .QN());
   DFF_X1 \buffer_reg[10][0][0][12]  (.D(\input_filter[0][0] [12]), .CK(n_56_7), 
      .Q(\buffer[10][0][0] [12]), .QN());
   DFF_X1 \buffer_reg[10][0][0][11]  (.D(\input_filter[0][0] [11]), .CK(n_56_7), 
      .Q(\buffer[10][0][0] [11]), .QN());
   DFF_X1 \buffer_reg[10][0][0][10]  (.D(\input_filter[0][0] [10]), .CK(n_56_7), 
      .Q(\buffer[10][0][0] [10]), .QN());
   DFF_X1 \buffer_reg[10][0][0][9]  (.D(\input_filter[0][0] [9]), .CK(n_56_7), 
      .Q(\buffer[10][0][0] [9]), .QN());
   DFF_X1 \buffer_reg[10][0][0][8]  (.D(\input_filter[0][0] [8]), .CK(n_56_7), 
      .Q(\buffer[10][0][0] [8]), .QN());
   DFF_X1 \buffer_reg[10][0][0][7]  (.D(\input_filter[0][0] [7]), .CK(n_56_7), 
      .Q(\buffer[10][0][0] [7]), .QN());
   DFF_X1 \buffer_reg[10][0][0][6]  (.D(\input_filter[0][0] [6]), .CK(n_56_7), 
      .Q(\buffer[10][0][0] [6]), .QN());
   DFF_X1 \buffer_reg[10][0][0][5]  (.D(\input_filter[0][0] [5]), .CK(n_56_7), 
      .Q(\buffer[10][0][0] [5]), .QN());
   DFF_X1 \buffer_reg[10][0][0][4]  (.D(\input_filter[0][0] [4]), .CK(n_56_7), 
      .Q(\buffer[10][0][0] [4]), .QN());
   DFF_X1 \buffer_reg[10][0][0][3]  (.D(\input_filter[0][0] [3]), .CK(n_56_7), 
      .Q(\buffer[10][0][0] [3]), .QN());
   DFF_X1 \buffer_reg[10][0][0][2]  (.D(\input_filter[0][0] [2]), .CK(n_56_7), 
      .Q(\buffer[10][0][0] [2]), .QN());
   DFF_X1 \buffer_reg[10][0][0][1]  (.D(\input_filter[0][0] [1]), .CK(n_56_7), 
      .Q(\buffer[10][0][0] [1]), .QN());
   DFF_X1 \buffer_reg[10][0][0][0]  (.D(\input_filter[0][0] [0]), .CK(n_56_7), 
      .Q(\buffer[10][0][0] [0]), .QN());
   DFF_X1 \buffer_reg[11][0][0][15]  (.D(\input_filter[0][0] [15]), .CK(n_56_8), 
      .Q(\buffer[11][0][0] [15]), .QN());
   DFF_X1 \buffer_reg[11][0][0][14]  (.D(\input_filter[0][0] [14]), .CK(n_56_8), 
      .Q(\buffer[11][0][0] [14]), .QN());
   DFF_X1 \buffer_reg[11][0][0][13]  (.D(\input_filter[0][0] [13]), .CK(n_56_8), 
      .Q(\buffer[11][0][0] [13]), .QN());
   DFF_X1 \buffer_reg[11][0][0][12]  (.D(\input_filter[0][0] [12]), .CK(n_56_8), 
      .Q(\buffer[11][0][0] [12]), .QN());
   DFF_X1 \buffer_reg[11][0][0][11]  (.D(\input_filter[0][0] [11]), .CK(n_56_8), 
      .Q(\buffer[11][0][0] [11]), .QN());
   DFF_X1 \buffer_reg[11][0][0][10]  (.D(\input_filter[0][0] [10]), .CK(n_56_8), 
      .Q(\buffer[11][0][0] [10]), .QN());
   DFF_X1 \buffer_reg[11][0][0][9]  (.D(\input_filter[0][0] [9]), .CK(n_56_8), 
      .Q(\buffer[11][0][0] [9]), .QN());
   DFF_X1 \buffer_reg[11][0][0][8]  (.D(\input_filter[0][0] [8]), .CK(n_56_8), 
      .Q(\buffer[11][0][0] [8]), .QN());
   DFF_X1 \buffer_reg[11][0][0][7]  (.D(\input_filter[0][0] [7]), .CK(n_56_8), 
      .Q(\buffer[11][0][0] [7]), .QN());
   DFF_X1 \buffer_reg[11][0][0][6]  (.D(\input_filter[0][0] [6]), .CK(n_56_8), 
      .Q(\buffer[11][0][0] [6]), .QN());
   DFF_X1 \buffer_reg[11][0][0][5]  (.D(\input_filter[0][0] [5]), .CK(n_56_8), 
      .Q(\buffer[11][0][0] [5]), .QN());
   DFF_X1 \buffer_reg[11][0][0][4]  (.D(\input_filter[0][0] [4]), .CK(n_56_8), 
      .Q(\buffer[11][0][0] [4]), .QN());
   DFF_X1 \buffer_reg[11][0][0][3]  (.D(\input_filter[0][0] [3]), .CK(n_56_8), 
      .Q(\buffer[11][0][0] [3]), .QN());
   DFF_X1 \buffer_reg[11][0][0][2]  (.D(\input_filter[0][0] [2]), .CK(n_56_8), 
      .Q(\buffer[11][0][0] [2]), .QN());
   DFF_X1 \buffer_reg[11][0][0][1]  (.D(\input_filter[0][0] [1]), .CK(n_56_8), 
      .Q(\buffer[11][0][0] [1]), .QN());
   DFF_X1 \buffer_reg[11][0][0][0]  (.D(\input_filter[0][0] [0]), .CK(n_56_8), 
      .Q(\buffer[11][0][0] [0]), .QN());
   DFF_X1 \buffer_reg[12][0][0][15]  (.D(\input_filter[0][0] [15]), .CK(n_56_9), 
      .Q(\buffer[12][0][0] [15]), .QN());
   DFF_X1 \buffer_reg[12][0][0][14]  (.D(\input_filter[0][0] [14]), .CK(n_56_9), 
      .Q(\buffer[12][0][0] [14]), .QN());
   DFF_X1 \buffer_reg[12][0][0][13]  (.D(\input_filter[0][0] [13]), .CK(n_56_9), 
      .Q(\buffer[12][0][0] [13]), .QN());
   DFF_X1 \buffer_reg[12][0][0][12]  (.D(\input_filter[0][0] [12]), .CK(n_56_9), 
      .Q(\buffer[12][0][0] [12]), .QN());
   DFF_X1 \buffer_reg[12][0][0][11]  (.D(\input_filter[0][0] [11]), .CK(n_56_9), 
      .Q(\buffer[12][0][0] [11]), .QN());
   DFF_X1 \buffer_reg[12][0][0][10]  (.D(\input_filter[0][0] [10]), .CK(n_56_9), 
      .Q(\buffer[12][0][0] [10]), .QN());
   DFF_X1 \buffer_reg[12][0][0][9]  (.D(\input_filter[0][0] [9]), .CK(n_56_9), 
      .Q(\buffer[12][0][0] [9]), .QN());
   DFF_X1 \buffer_reg[12][0][0][8]  (.D(\input_filter[0][0] [8]), .CK(n_56_9), 
      .Q(\buffer[12][0][0] [8]), .QN());
   DFF_X1 \buffer_reg[12][0][0][7]  (.D(\input_filter[0][0] [7]), .CK(n_56_9), 
      .Q(\buffer[12][0][0] [7]), .QN());
   DFF_X1 \buffer_reg[12][0][0][6]  (.D(\input_filter[0][0] [6]), .CK(n_56_9), 
      .Q(\buffer[12][0][0] [6]), .QN());
   DFF_X1 \buffer_reg[12][0][0][5]  (.D(\input_filter[0][0] [5]), .CK(n_56_9), 
      .Q(\buffer[12][0][0] [5]), .QN());
   DFF_X1 \buffer_reg[12][0][0][4]  (.D(\input_filter[0][0] [4]), .CK(n_56_9), 
      .Q(\buffer[12][0][0] [4]), .QN());
   DFF_X1 \buffer_reg[12][0][0][3]  (.D(\input_filter[0][0] [3]), .CK(n_56_9), 
      .Q(\buffer[12][0][0] [3]), .QN());
   DFF_X1 \buffer_reg[12][0][0][2]  (.D(\input_filter[0][0] [2]), .CK(n_56_9), 
      .Q(\buffer[12][0][0] [2]), .QN());
   DFF_X1 \buffer_reg[12][0][0][1]  (.D(\input_filter[0][0] [1]), .CK(n_56_9), 
      .Q(\buffer[12][0][0] [1]), .QN());
   DFF_X1 \buffer_reg[12][0][0][0]  (.D(\input_filter[0][0] [0]), .CK(n_56_9), 
      .Q(\buffer[12][0][0] [0]), .QN());
   DFF_X1 \buffer_reg[13][0][0][15]  (.D(\input_filter[0][0] [15]), .CK(n_56_10), 
      .Q(\buffer[13][0][0] [15]), .QN());
   DFF_X1 \buffer_reg[13][0][0][14]  (.D(\input_filter[0][0] [14]), .CK(n_56_10), 
      .Q(\buffer[13][0][0] [14]), .QN());
   DFF_X1 \buffer_reg[13][0][0][13]  (.D(\input_filter[0][0] [13]), .CK(n_56_10), 
      .Q(\buffer[13][0][0] [13]), .QN());
   DFF_X1 \buffer_reg[13][0][0][12]  (.D(\input_filter[0][0] [12]), .CK(n_56_10), 
      .Q(\buffer[13][0][0] [12]), .QN());
   DFF_X1 \buffer_reg[13][0][0][11]  (.D(\input_filter[0][0] [11]), .CK(n_56_10), 
      .Q(\buffer[13][0][0] [11]), .QN());
   DFF_X1 \buffer_reg[13][0][0][10]  (.D(\input_filter[0][0] [10]), .CK(n_56_10), 
      .Q(\buffer[13][0][0] [10]), .QN());
   DFF_X1 \buffer_reg[13][0][0][9]  (.D(\input_filter[0][0] [9]), .CK(n_56_10), 
      .Q(\buffer[13][0][0] [9]), .QN());
   DFF_X1 \buffer_reg[13][0][0][8]  (.D(\input_filter[0][0] [8]), .CK(n_56_10), 
      .Q(\buffer[13][0][0] [8]), .QN());
   DFF_X1 \buffer_reg[13][0][0][7]  (.D(\input_filter[0][0] [7]), .CK(n_56_10), 
      .Q(\buffer[13][0][0] [7]), .QN());
   DFF_X1 \buffer_reg[13][0][0][6]  (.D(\input_filter[0][0] [6]), .CK(n_56_10), 
      .Q(\buffer[13][0][0] [6]), .QN());
   DFF_X1 \buffer_reg[13][0][0][5]  (.D(\input_filter[0][0] [5]), .CK(n_56_10), 
      .Q(\buffer[13][0][0] [5]), .QN());
   DFF_X1 \buffer_reg[13][0][0][4]  (.D(\input_filter[0][0] [4]), .CK(n_56_10), 
      .Q(\buffer[13][0][0] [4]), .QN());
   DFF_X1 \buffer_reg[13][0][0][3]  (.D(\input_filter[0][0] [3]), .CK(n_56_10), 
      .Q(\buffer[13][0][0] [3]), .QN());
   DFF_X1 \buffer_reg[13][0][0][2]  (.D(\input_filter[0][0] [2]), .CK(n_56_10), 
      .Q(\buffer[13][0][0] [2]), .QN());
   DFF_X1 \buffer_reg[13][0][0][1]  (.D(\input_filter[0][0] [1]), .CK(n_56_10), 
      .Q(\buffer[13][0][0] [1]), .QN());
   DFF_X1 \buffer_reg[13][0][0][0]  (.D(\input_filter[0][0] [0]), .CK(n_56_10), 
      .Q(\buffer[13][0][0] [0]), .QN());
   DFF_X1 \buffer_reg[14][0][0][15]  (.D(\input_filter[0][0] [15]), .CK(n_56_11), 
      .Q(\buffer[14][0][0] [15]), .QN());
   DFF_X1 \buffer_reg[14][0][0][14]  (.D(\input_filter[0][0] [14]), .CK(n_56_11), 
      .Q(\buffer[14][0][0] [14]), .QN());
   DFF_X1 \buffer_reg[14][0][0][13]  (.D(\input_filter[0][0] [13]), .CK(n_56_11), 
      .Q(\buffer[14][0][0] [13]), .QN());
   DFF_X1 \buffer_reg[14][0][0][12]  (.D(\input_filter[0][0] [12]), .CK(n_56_11), 
      .Q(\buffer[14][0][0] [12]), .QN());
   DFF_X1 \buffer_reg[14][0][0][11]  (.D(\input_filter[0][0] [11]), .CK(n_56_11), 
      .Q(\buffer[14][0][0] [11]), .QN());
   DFF_X1 \buffer_reg[14][0][0][10]  (.D(\input_filter[0][0] [10]), .CK(n_56_11), 
      .Q(\buffer[14][0][0] [10]), .QN());
   DFF_X1 \buffer_reg[14][0][0][9]  (.D(\input_filter[0][0] [9]), .CK(n_56_11), 
      .Q(\buffer[14][0][0] [9]), .QN());
   DFF_X1 \buffer_reg[14][0][0][8]  (.D(\input_filter[0][0] [8]), .CK(n_56_11), 
      .Q(\buffer[14][0][0] [8]), .QN());
   DFF_X1 \buffer_reg[14][0][0][7]  (.D(\input_filter[0][0] [7]), .CK(n_56_11), 
      .Q(\buffer[14][0][0] [7]), .QN());
   DFF_X1 \buffer_reg[14][0][0][6]  (.D(\input_filter[0][0] [6]), .CK(n_56_11), 
      .Q(\buffer[14][0][0] [6]), .QN());
   DFF_X1 \buffer_reg[14][0][0][5]  (.D(\input_filter[0][0] [5]), .CK(n_56_11), 
      .Q(\buffer[14][0][0] [5]), .QN());
   DFF_X1 \buffer_reg[14][0][0][4]  (.D(\input_filter[0][0] [4]), .CK(n_56_11), 
      .Q(\buffer[14][0][0] [4]), .QN());
   DFF_X1 \buffer_reg[14][0][0][3]  (.D(\input_filter[0][0] [3]), .CK(n_56_11), 
      .Q(\buffer[14][0][0] [3]), .QN());
   DFF_X1 \buffer_reg[14][0][0][2]  (.D(\input_filter[0][0] [2]), .CK(n_56_11), 
      .Q(\buffer[14][0][0] [2]), .QN());
   DFF_X1 \buffer_reg[14][0][0][1]  (.D(\input_filter[0][0] [1]), .CK(n_56_11), 
      .Q(\buffer[14][0][0] [1]), .QN());
   DFF_X1 \buffer_reg[14][0][0][0]  (.D(\input_filter[0][0] [0]), .CK(n_56_11), 
      .Q(\buffer[14][0][0] [0]), .QN());
   DFF_X1 \buffer_reg[0][0][1][15]  (.D(\input_filter[0][1] [15]), .CK(n_56_12), 
      .Q(\buffer[0][0][1] [15]), .QN());
   DFF_X1 \buffer_reg[0][0][1][14]  (.D(\input_filter[0][1] [14]), .CK(n_56_12), 
      .Q(\buffer[0][0][1] [14]), .QN());
   DFF_X1 \buffer_reg[0][0][1][13]  (.D(\input_filter[0][1] [13]), .CK(n_56_12), 
      .Q(\buffer[0][0][1] [13]), .QN());
   DFF_X1 \buffer_reg[0][0][1][12]  (.D(\input_filter[0][1] [12]), .CK(n_56_12), 
      .Q(\buffer[0][0][1] [12]), .QN());
   DFF_X1 \buffer_reg[0][0][1][11]  (.D(\input_filter[0][1] [11]), .CK(n_56_12), 
      .Q(\buffer[0][0][1] [11]), .QN());
   DFF_X1 \buffer_reg[0][0][1][10]  (.D(\input_filter[0][1] [10]), .CK(n_56_12), 
      .Q(\buffer[0][0][1] [10]), .QN());
   DFF_X1 \buffer_reg[0][0][1][9]  (.D(\input_filter[0][1] [9]), .CK(n_56_12), 
      .Q(\buffer[0][0][1] [9]), .QN());
   DFF_X1 \buffer_reg[0][0][1][8]  (.D(\input_filter[0][1] [8]), .CK(n_56_12), 
      .Q(\buffer[0][0][1] [8]), .QN());
   DFF_X1 \buffer_reg[0][0][1][7]  (.D(\input_filter[0][1] [7]), .CK(n_56_12), 
      .Q(\buffer[0][0][1] [7]), .QN());
   DFF_X1 \buffer_reg[0][0][1][6]  (.D(\input_filter[0][1] [6]), .CK(n_56_12), 
      .Q(\buffer[0][0][1] [6]), .QN());
   DFF_X1 \buffer_reg[0][0][1][5]  (.D(\input_filter[0][1] [5]), .CK(n_56_12), 
      .Q(\buffer[0][0][1] [5]), .QN());
   DFF_X1 \buffer_reg[0][0][1][4]  (.D(\input_filter[0][1] [4]), .CK(n_56_12), 
      .Q(\buffer[0][0][1] [4]), .QN());
   DFF_X1 \buffer_reg[0][0][1][3]  (.D(\input_filter[0][1] [3]), .CK(n_56_12), 
      .Q(\buffer[0][0][1] [3]), .QN());
   DFF_X1 \buffer_reg[0][0][1][2]  (.D(\input_filter[0][1] [2]), .CK(n_56_12), 
      .Q(\buffer[0][0][1] [2]), .QN());
   DFF_X1 \buffer_reg[0][0][1][1]  (.D(\input_filter[0][1] [1]), .CK(n_56_12), 
      .Q(\buffer[0][0][1] [1]), .QN());
   DFF_X1 \buffer_reg[0][0][1][0]  (.D(\input_filter[0][1] [0]), .CK(n_56_12), 
      .Q(\buffer[0][0][1] [0]), .QN());
   DFF_X1 \buffer_reg[1][0][1][15]  (.D(\input_filter[0][1] [15]), .CK(n_56_13), 
      .Q(\buffer[1][0][1] [15]), .QN());
   DFF_X1 \buffer_reg[1][0][1][14]  (.D(\input_filter[0][1] [14]), .CK(n_56_13), 
      .Q(\buffer[1][0][1] [14]), .QN());
   DFF_X1 \buffer_reg[1][0][1][13]  (.D(\input_filter[0][1] [13]), .CK(n_56_13), 
      .Q(\buffer[1][0][1] [13]), .QN());
   DFF_X1 \buffer_reg[1][0][1][12]  (.D(\input_filter[0][1] [12]), .CK(n_56_13), 
      .Q(\buffer[1][0][1] [12]), .QN());
   DFF_X1 \buffer_reg[1][0][1][11]  (.D(\input_filter[0][1] [11]), .CK(n_56_13), 
      .Q(\buffer[1][0][1] [11]), .QN());
   DFF_X1 \buffer_reg[1][0][1][10]  (.D(\input_filter[0][1] [10]), .CK(n_56_13), 
      .Q(\buffer[1][0][1] [10]), .QN());
   DFF_X1 \buffer_reg[1][0][1][9]  (.D(\input_filter[0][1] [9]), .CK(n_56_13), 
      .Q(\buffer[1][0][1] [9]), .QN());
   DFF_X1 \buffer_reg[1][0][1][8]  (.D(\input_filter[0][1] [8]), .CK(n_56_13), 
      .Q(\buffer[1][0][1] [8]), .QN());
   DFF_X1 \buffer_reg[1][0][1][7]  (.D(\input_filter[0][1] [7]), .CK(n_56_13), 
      .Q(\buffer[1][0][1] [7]), .QN());
   DFF_X1 \buffer_reg[1][0][1][6]  (.D(\input_filter[0][1] [6]), .CK(n_56_13), 
      .Q(\buffer[1][0][1] [6]), .QN());
   DFF_X1 \buffer_reg[1][0][1][5]  (.D(\input_filter[0][1] [5]), .CK(n_56_13), 
      .Q(\buffer[1][0][1] [5]), .QN());
   DFF_X1 \buffer_reg[1][0][1][4]  (.D(\input_filter[0][1] [4]), .CK(n_56_13), 
      .Q(\buffer[1][0][1] [4]), .QN());
   DFF_X1 \buffer_reg[1][0][1][3]  (.D(\input_filter[0][1] [3]), .CK(n_56_13), 
      .Q(\buffer[1][0][1] [3]), .QN());
   DFF_X1 \buffer_reg[1][0][1][2]  (.D(\input_filter[0][1] [2]), .CK(n_56_13), 
      .Q(\buffer[1][0][1] [2]), .QN());
   DFF_X1 \buffer_reg[1][0][1][1]  (.D(\input_filter[0][1] [1]), .CK(n_56_13), 
      .Q(\buffer[1][0][1] [1]), .QN());
   DFF_X1 \buffer_reg[1][0][1][0]  (.D(\input_filter[0][1] [0]), .CK(n_56_13), 
      .Q(\buffer[1][0][1] [0]), .QN());
   DFF_X1 \buffer_reg[2][0][1][15]  (.D(\input_filter[0][1] [15]), .CK(n_56_14), 
      .Q(\buffer[2][0][1] [15]), .QN());
   DFF_X1 \buffer_reg[2][0][1][14]  (.D(\input_filter[0][1] [14]), .CK(n_56_14), 
      .Q(\buffer[2][0][1] [14]), .QN());
   DFF_X1 \buffer_reg[2][0][1][13]  (.D(\input_filter[0][1] [13]), .CK(n_56_14), 
      .Q(\buffer[2][0][1] [13]), .QN());
   DFF_X1 \buffer_reg[2][0][1][12]  (.D(\input_filter[0][1] [12]), .CK(n_56_14), 
      .Q(\buffer[2][0][1] [12]), .QN());
   DFF_X1 \buffer_reg[2][0][1][11]  (.D(\input_filter[0][1] [11]), .CK(n_56_14), 
      .Q(\buffer[2][0][1] [11]), .QN());
   DFF_X1 \buffer_reg[2][0][1][10]  (.D(\input_filter[0][1] [10]), .CK(n_56_14), 
      .Q(\buffer[2][0][1] [10]), .QN());
   DFF_X1 \buffer_reg[2][0][1][9]  (.D(\input_filter[0][1] [9]), .CK(n_56_14), 
      .Q(\buffer[2][0][1] [9]), .QN());
   DFF_X1 \buffer_reg[2][0][1][8]  (.D(\input_filter[0][1] [8]), .CK(n_56_14), 
      .Q(\buffer[2][0][1] [8]), .QN());
   DFF_X1 \buffer_reg[2][0][1][7]  (.D(\input_filter[0][1] [7]), .CK(n_56_14), 
      .Q(\buffer[2][0][1] [7]), .QN());
   DFF_X1 \buffer_reg[2][0][1][6]  (.D(\input_filter[0][1] [6]), .CK(n_56_14), 
      .Q(\buffer[2][0][1] [6]), .QN());
   DFF_X1 \buffer_reg[2][0][1][5]  (.D(\input_filter[0][1] [5]), .CK(n_56_14), 
      .Q(\buffer[2][0][1] [5]), .QN());
   DFF_X1 \buffer_reg[2][0][1][4]  (.D(\input_filter[0][1] [4]), .CK(n_56_14), 
      .Q(\buffer[2][0][1] [4]), .QN());
   DFF_X1 \buffer_reg[2][0][1][3]  (.D(\input_filter[0][1] [3]), .CK(n_56_14), 
      .Q(\buffer[2][0][1] [3]), .QN());
   DFF_X1 \buffer_reg[2][0][1][2]  (.D(\input_filter[0][1] [2]), .CK(n_56_14), 
      .Q(\buffer[2][0][1] [2]), .QN());
   DFF_X1 \buffer_reg[2][0][1][1]  (.D(\input_filter[0][1] [1]), .CK(n_56_14), 
      .Q(\buffer[2][0][1] [1]), .QN());
   DFF_X1 \buffer_reg[2][0][1][0]  (.D(\input_filter[0][1] [0]), .CK(n_56_14), 
      .Q(\buffer[2][0][1] [0]), .QN());
   DFF_X1 \buffer_reg[3][0][1][15]  (.D(\input_filter[0][1] [15]), .CK(n_56_0), 
      .Q(\buffer[3][0][1] [15]), .QN());
   DFF_X1 \buffer_reg[3][0][1][14]  (.D(\input_filter[0][1] [14]), .CK(n_56_0), 
      .Q(\buffer[3][0][1] [14]), .QN());
   DFF_X1 \buffer_reg[3][0][1][13]  (.D(\input_filter[0][1] [13]), .CK(n_56_0), 
      .Q(\buffer[3][0][1] [13]), .QN());
   DFF_X1 \buffer_reg[3][0][1][12]  (.D(\input_filter[0][1] [12]), .CK(n_56_0), 
      .Q(\buffer[3][0][1] [12]), .QN());
   DFF_X1 \buffer_reg[3][0][1][11]  (.D(\input_filter[0][1] [11]), .CK(n_56_0), 
      .Q(\buffer[3][0][1] [11]), .QN());
   DFF_X1 \buffer_reg[3][0][1][10]  (.D(\input_filter[0][1] [10]), .CK(n_56_0), 
      .Q(\buffer[3][0][1] [10]), .QN());
   DFF_X1 \buffer_reg[3][0][1][9]  (.D(\input_filter[0][1] [9]), .CK(n_56_0), 
      .Q(\buffer[3][0][1] [9]), .QN());
   DFF_X1 \buffer_reg[3][0][1][8]  (.D(\input_filter[0][1] [8]), .CK(n_56_0), 
      .Q(\buffer[3][0][1] [8]), .QN());
   DFF_X1 \buffer_reg[3][0][1][7]  (.D(\input_filter[0][1] [7]), .CK(n_56_0), 
      .Q(\buffer[3][0][1] [7]), .QN());
   DFF_X1 \buffer_reg[3][0][1][6]  (.D(\input_filter[0][1] [6]), .CK(n_56_0), 
      .Q(\buffer[3][0][1] [6]), .QN());
   DFF_X1 \buffer_reg[3][0][1][5]  (.D(\input_filter[0][1] [5]), .CK(n_56_0), 
      .Q(\buffer[3][0][1] [5]), .QN());
   DFF_X1 \buffer_reg[3][0][1][4]  (.D(\input_filter[0][1] [4]), .CK(n_56_0), 
      .Q(\buffer[3][0][1] [4]), .QN());
   DFF_X1 \buffer_reg[3][0][1][3]  (.D(\input_filter[0][1] [3]), .CK(n_56_0), 
      .Q(\buffer[3][0][1] [3]), .QN());
   DFF_X1 \buffer_reg[3][0][1][2]  (.D(\input_filter[0][1] [2]), .CK(n_56_0), 
      .Q(\buffer[3][0][1] [2]), .QN());
   DFF_X1 \buffer_reg[3][0][1][1]  (.D(\input_filter[0][1] [1]), .CK(n_56_0), 
      .Q(\buffer[3][0][1] [1]), .QN());
   DFF_X1 \buffer_reg[3][0][1][0]  (.D(\input_filter[0][1] [0]), .CK(n_56_0), 
      .Q(\buffer[3][0][1] [0]), .QN());
   DFF_X1 \buffer_reg[4][0][1][15]  (.D(\input_filter[0][1] [15]), .CK(n_56_1), 
      .Q(\buffer[4][0][1] [15]), .QN());
   DFF_X1 \buffer_reg[4][0][1][14]  (.D(\input_filter[0][1] [14]), .CK(n_56_1), 
      .Q(\buffer[4][0][1] [14]), .QN());
   DFF_X1 \buffer_reg[4][0][1][13]  (.D(\input_filter[0][1] [13]), .CK(n_56_1), 
      .Q(\buffer[4][0][1] [13]), .QN());
   DFF_X1 \buffer_reg[4][0][1][12]  (.D(\input_filter[0][1] [12]), .CK(n_56_1), 
      .Q(\buffer[4][0][1] [12]), .QN());
   DFF_X1 \buffer_reg[4][0][1][11]  (.D(\input_filter[0][1] [11]), .CK(n_56_1), 
      .Q(\buffer[4][0][1] [11]), .QN());
   DFF_X1 \buffer_reg[4][0][1][10]  (.D(\input_filter[0][1] [10]), .CK(n_56_1), 
      .Q(\buffer[4][0][1] [10]), .QN());
   DFF_X1 \buffer_reg[4][0][1][9]  (.D(\input_filter[0][1] [9]), .CK(n_56_1), 
      .Q(\buffer[4][0][1] [9]), .QN());
   DFF_X1 \buffer_reg[4][0][1][8]  (.D(\input_filter[0][1] [8]), .CK(n_56_1), 
      .Q(\buffer[4][0][1] [8]), .QN());
   DFF_X1 \buffer_reg[4][0][1][7]  (.D(\input_filter[0][1] [7]), .CK(n_56_1), 
      .Q(\buffer[4][0][1] [7]), .QN());
   DFF_X1 \buffer_reg[4][0][1][6]  (.D(\input_filter[0][1] [6]), .CK(n_56_1), 
      .Q(\buffer[4][0][1] [6]), .QN());
   DFF_X1 \buffer_reg[4][0][1][5]  (.D(\input_filter[0][1] [5]), .CK(n_56_1), 
      .Q(\buffer[4][0][1] [5]), .QN());
   DFF_X1 \buffer_reg[4][0][1][4]  (.D(\input_filter[0][1] [4]), .CK(n_56_1), 
      .Q(\buffer[4][0][1] [4]), .QN());
   DFF_X1 \buffer_reg[4][0][1][3]  (.D(\input_filter[0][1] [3]), .CK(n_56_1), 
      .Q(\buffer[4][0][1] [3]), .QN());
   DFF_X1 \buffer_reg[4][0][1][2]  (.D(\input_filter[0][1] [2]), .CK(n_56_1), 
      .Q(\buffer[4][0][1] [2]), .QN());
   DFF_X1 \buffer_reg[4][0][1][1]  (.D(\input_filter[0][1] [1]), .CK(n_56_1), 
      .Q(\buffer[4][0][1] [1]), .QN());
   DFF_X1 \buffer_reg[4][0][1][0]  (.D(\input_filter[0][1] [0]), .CK(n_56_1), 
      .Q(\buffer[4][0][1] [0]), .QN());
   DFF_X1 \buffer_reg[5][0][1][15]  (.D(\input_filter[0][1] [15]), .CK(n_56_2), 
      .Q(\buffer[5][0][1] [15]), .QN());
   DFF_X1 \buffer_reg[5][0][1][14]  (.D(\input_filter[0][1] [14]), .CK(n_56_2), 
      .Q(\buffer[5][0][1] [14]), .QN());
   DFF_X1 \buffer_reg[5][0][1][13]  (.D(\input_filter[0][1] [13]), .CK(n_56_2), 
      .Q(\buffer[5][0][1] [13]), .QN());
   DFF_X1 \buffer_reg[5][0][1][12]  (.D(\input_filter[0][1] [12]), .CK(n_56_2), 
      .Q(\buffer[5][0][1] [12]), .QN());
   DFF_X1 \buffer_reg[5][0][1][11]  (.D(\input_filter[0][1] [11]), .CK(n_56_2), 
      .Q(\buffer[5][0][1] [11]), .QN());
   DFF_X1 \buffer_reg[5][0][1][10]  (.D(\input_filter[0][1] [10]), .CK(n_56_2), 
      .Q(\buffer[5][0][1] [10]), .QN());
   DFF_X1 \buffer_reg[5][0][1][9]  (.D(\input_filter[0][1] [9]), .CK(n_56_2), 
      .Q(\buffer[5][0][1] [9]), .QN());
   DFF_X1 \buffer_reg[5][0][1][8]  (.D(\input_filter[0][1] [8]), .CK(n_56_2), 
      .Q(\buffer[5][0][1] [8]), .QN());
   DFF_X1 \buffer_reg[5][0][1][7]  (.D(\input_filter[0][1] [7]), .CK(n_56_2), 
      .Q(\buffer[5][0][1] [7]), .QN());
   DFF_X1 \buffer_reg[5][0][1][6]  (.D(\input_filter[0][1] [6]), .CK(n_56_2), 
      .Q(\buffer[5][0][1] [6]), .QN());
   DFF_X1 \buffer_reg[5][0][1][5]  (.D(\input_filter[0][1] [5]), .CK(n_56_2), 
      .Q(\buffer[5][0][1] [5]), .QN());
   DFF_X1 \buffer_reg[5][0][1][4]  (.D(\input_filter[0][1] [4]), .CK(n_56_2), 
      .Q(\buffer[5][0][1] [4]), .QN());
   DFF_X1 \buffer_reg[5][0][1][3]  (.D(\input_filter[0][1] [3]), .CK(n_56_2), 
      .Q(\buffer[5][0][1] [3]), .QN());
   DFF_X1 \buffer_reg[5][0][1][2]  (.D(\input_filter[0][1] [2]), .CK(n_56_2), 
      .Q(\buffer[5][0][1] [2]), .QN());
   DFF_X1 \buffer_reg[5][0][1][1]  (.D(\input_filter[0][1] [1]), .CK(n_56_2), 
      .Q(\buffer[5][0][1] [1]), .QN());
   DFF_X1 \buffer_reg[5][0][1][0]  (.D(\input_filter[0][1] [0]), .CK(n_56_2), 
      .Q(\buffer[5][0][1] [0]), .QN());
   DFF_X1 \buffer_reg[6][0][1][15]  (.D(\input_filter[0][1] [15]), .CK(n_56_3), 
      .Q(\buffer[6][0][1] [15]), .QN());
   DFF_X1 \buffer_reg[6][0][1][14]  (.D(\input_filter[0][1] [14]), .CK(n_56_3), 
      .Q(\buffer[6][0][1] [14]), .QN());
   DFF_X1 \buffer_reg[6][0][1][13]  (.D(\input_filter[0][1] [13]), .CK(n_56_3), 
      .Q(\buffer[6][0][1] [13]), .QN());
   DFF_X1 \buffer_reg[6][0][1][12]  (.D(\input_filter[0][1] [12]), .CK(n_56_3), 
      .Q(\buffer[6][0][1] [12]), .QN());
   DFF_X1 \buffer_reg[6][0][1][11]  (.D(\input_filter[0][1] [11]), .CK(n_56_3), 
      .Q(\buffer[6][0][1] [11]), .QN());
   DFF_X1 \buffer_reg[6][0][1][10]  (.D(\input_filter[0][1] [10]), .CK(n_56_3), 
      .Q(\buffer[6][0][1] [10]), .QN());
   DFF_X1 \buffer_reg[6][0][1][9]  (.D(\input_filter[0][1] [9]), .CK(n_56_3), 
      .Q(\buffer[6][0][1] [9]), .QN());
   DFF_X1 \buffer_reg[6][0][1][8]  (.D(\input_filter[0][1] [8]), .CK(n_56_3), 
      .Q(\buffer[6][0][1] [8]), .QN());
   DFF_X1 \buffer_reg[6][0][1][7]  (.D(\input_filter[0][1] [7]), .CK(n_56_3), 
      .Q(\buffer[6][0][1] [7]), .QN());
   DFF_X1 \buffer_reg[6][0][1][6]  (.D(\input_filter[0][1] [6]), .CK(n_56_3), 
      .Q(\buffer[6][0][1] [6]), .QN());
   DFF_X1 \buffer_reg[6][0][1][5]  (.D(\input_filter[0][1] [5]), .CK(n_56_3), 
      .Q(\buffer[6][0][1] [5]), .QN());
   DFF_X1 \buffer_reg[6][0][1][4]  (.D(\input_filter[0][1] [4]), .CK(n_56_3), 
      .Q(\buffer[6][0][1] [4]), .QN());
   DFF_X1 \buffer_reg[6][0][1][3]  (.D(\input_filter[0][1] [3]), .CK(n_56_3), 
      .Q(\buffer[6][0][1] [3]), .QN());
   DFF_X1 \buffer_reg[6][0][1][2]  (.D(\input_filter[0][1] [2]), .CK(n_56_3), 
      .Q(\buffer[6][0][1] [2]), .QN());
   DFF_X1 \buffer_reg[6][0][1][1]  (.D(\input_filter[0][1] [1]), .CK(n_56_3), 
      .Q(\buffer[6][0][1] [1]), .QN());
   DFF_X1 \buffer_reg[6][0][1][0]  (.D(\input_filter[0][1] [0]), .CK(n_56_3), 
      .Q(\buffer[6][0][1] [0]), .QN());
   DFF_X1 \buffer_reg[7][0][1][15]  (.D(\input_filter[0][1] [15]), .CK(n_56_4), 
      .Q(\buffer[7][0][1] [15]), .QN());
   DFF_X1 \buffer_reg[7][0][1][14]  (.D(\input_filter[0][1] [14]), .CK(n_56_4), 
      .Q(\buffer[7][0][1] [14]), .QN());
   DFF_X1 \buffer_reg[7][0][1][13]  (.D(\input_filter[0][1] [13]), .CK(n_56_4), 
      .Q(\buffer[7][0][1] [13]), .QN());
   DFF_X1 \buffer_reg[7][0][1][12]  (.D(\input_filter[0][1] [12]), .CK(n_56_4), 
      .Q(\buffer[7][0][1] [12]), .QN());
   DFF_X1 \buffer_reg[7][0][1][11]  (.D(\input_filter[0][1] [11]), .CK(n_56_4), 
      .Q(\buffer[7][0][1] [11]), .QN());
   DFF_X1 \buffer_reg[7][0][1][10]  (.D(\input_filter[0][1] [10]), .CK(n_56_4), 
      .Q(\buffer[7][0][1] [10]), .QN());
   DFF_X1 \buffer_reg[7][0][1][9]  (.D(\input_filter[0][1] [9]), .CK(n_56_4), 
      .Q(\buffer[7][0][1] [9]), .QN());
   DFF_X1 \buffer_reg[7][0][1][8]  (.D(\input_filter[0][1] [8]), .CK(n_56_4), 
      .Q(\buffer[7][0][1] [8]), .QN());
   DFF_X1 \buffer_reg[7][0][1][7]  (.D(\input_filter[0][1] [7]), .CK(n_56_4), 
      .Q(\buffer[7][0][1] [7]), .QN());
   DFF_X1 \buffer_reg[7][0][1][6]  (.D(\input_filter[0][1] [6]), .CK(n_56_4), 
      .Q(\buffer[7][0][1] [6]), .QN());
   DFF_X1 \buffer_reg[7][0][1][5]  (.D(\input_filter[0][1] [5]), .CK(n_56_4), 
      .Q(\buffer[7][0][1] [5]), .QN());
   DFF_X1 \buffer_reg[7][0][1][4]  (.D(\input_filter[0][1] [4]), .CK(n_56_4), 
      .Q(\buffer[7][0][1] [4]), .QN());
   DFF_X1 \buffer_reg[7][0][1][3]  (.D(\input_filter[0][1] [3]), .CK(n_56_4), 
      .Q(\buffer[7][0][1] [3]), .QN());
   DFF_X1 \buffer_reg[7][0][1][2]  (.D(\input_filter[0][1] [2]), .CK(n_56_4), 
      .Q(\buffer[7][0][1] [2]), .QN());
   DFF_X1 \buffer_reg[7][0][1][1]  (.D(\input_filter[0][1] [1]), .CK(n_56_4), 
      .Q(\buffer[7][0][1] [1]), .QN());
   DFF_X1 \buffer_reg[7][0][1][0]  (.D(\input_filter[0][1] [0]), .CK(n_56_4), 
      .Q(\buffer[7][0][1] [0]), .QN());
   DFF_X1 \buffer_reg[8][0][1][15]  (.D(\input_filter[0][1] [15]), .CK(n_56_5), 
      .Q(\buffer[8][0][1] [15]), .QN());
   DFF_X1 \buffer_reg[8][0][1][14]  (.D(\input_filter[0][1] [14]), .CK(n_56_5), 
      .Q(\buffer[8][0][1] [14]), .QN());
   DFF_X1 \buffer_reg[8][0][1][13]  (.D(\input_filter[0][1] [13]), .CK(n_56_5), 
      .Q(\buffer[8][0][1] [13]), .QN());
   DFF_X1 \buffer_reg[8][0][1][12]  (.D(\input_filter[0][1] [12]), .CK(n_56_5), 
      .Q(\buffer[8][0][1] [12]), .QN());
   DFF_X1 \buffer_reg[8][0][1][11]  (.D(\input_filter[0][1] [11]), .CK(n_56_5), 
      .Q(\buffer[8][0][1] [11]), .QN());
   DFF_X1 \buffer_reg[8][0][1][10]  (.D(\input_filter[0][1] [10]), .CK(n_56_5), 
      .Q(\buffer[8][0][1] [10]), .QN());
   DFF_X1 \buffer_reg[8][0][1][9]  (.D(\input_filter[0][1] [9]), .CK(n_56_5), 
      .Q(\buffer[8][0][1] [9]), .QN());
   DFF_X1 \buffer_reg[8][0][1][8]  (.D(\input_filter[0][1] [8]), .CK(n_56_5), 
      .Q(\buffer[8][0][1] [8]), .QN());
   DFF_X1 \buffer_reg[8][0][1][7]  (.D(\input_filter[0][1] [7]), .CK(n_56_5), 
      .Q(\buffer[8][0][1] [7]), .QN());
   DFF_X1 \buffer_reg[8][0][1][6]  (.D(\input_filter[0][1] [6]), .CK(n_56_5), 
      .Q(\buffer[8][0][1] [6]), .QN());
   DFF_X1 \buffer_reg[8][0][1][5]  (.D(\input_filter[0][1] [5]), .CK(n_56_5), 
      .Q(\buffer[8][0][1] [5]), .QN());
   DFF_X1 \buffer_reg[8][0][1][4]  (.D(\input_filter[0][1] [4]), .CK(n_56_5), 
      .Q(\buffer[8][0][1] [4]), .QN());
   DFF_X1 \buffer_reg[8][0][1][3]  (.D(\input_filter[0][1] [3]), .CK(n_56_5), 
      .Q(\buffer[8][0][1] [3]), .QN());
   DFF_X1 \buffer_reg[8][0][1][2]  (.D(\input_filter[0][1] [2]), .CK(n_56_5), 
      .Q(\buffer[8][0][1] [2]), .QN());
   DFF_X1 \buffer_reg[8][0][1][1]  (.D(\input_filter[0][1] [1]), .CK(n_56_5), 
      .Q(\buffer[8][0][1] [1]), .QN());
   DFF_X1 \buffer_reg[8][0][1][0]  (.D(\input_filter[0][1] [0]), .CK(n_56_5), 
      .Q(\buffer[8][0][1] [0]), .QN());
   DFF_X1 \buffer_reg[9][0][1][15]  (.D(\input_filter[0][1] [15]), .CK(n_56_6), 
      .Q(\buffer[9][0][1] [15]), .QN());
   DFF_X1 \buffer_reg[9][0][1][14]  (.D(\input_filter[0][1] [14]), .CK(n_56_6), 
      .Q(\buffer[9][0][1] [14]), .QN());
   DFF_X1 \buffer_reg[9][0][1][13]  (.D(\input_filter[0][1] [13]), .CK(n_56_6), 
      .Q(\buffer[9][0][1] [13]), .QN());
   DFF_X1 \buffer_reg[9][0][1][12]  (.D(\input_filter[0][1] [12]), .CK(n_56_6), 
      .Q(\buffer[9][0][1] [12]), .QN());
   DFF_X1 \buffer_reg[9][0][1][11]  (.D(\input_filter[0][1] [11]), .CK(n_56_6), 
      .Q(\buffer[9][0][1] [11]), .QN());
   DFF_X1 \buffer_reg[9][0][1][10]  (.D(\input_filter[0][1] [10]), .CK(n_56_6), 
      .Q(\buffer[9][0][1] [10]), .QN());
   DFF_X1 \buffer_reg[9][0][1][9]  (.D(\input_filter[0][1] [9]), .CK(n_56_6), 
      .Q(\buffer[9][0][1] [9]), .QN());
   DFF_X1 \buffer_reg[9][0][1][8]  (.D(\input_filter[0][1] [8]), .CK(n_56_6), 
      .Q(\buffer[9][0][1] [8]), .QN());
   DFF_X1 \buffer_reg[9][0][1][7]  (.D(\input_filter[0][1] [7]), .CK(n_56_6), 
      .Q(\buffer[9][0][1] [7]), .QN());
   DFF_X1 \buffer_reg[9][0][1][6]  (.D(\input_filter[0][1] [6]), .CK(n_56_6), 
      .Q(\buffer[9][0][1] [6]), .QN());
   DFF_X1 \buffer_reg[9][0][1][5]  (.D(\input_filter[0][1] [5]), .CK(n_56_6), 
      .Q(\buffer[9][0][1] [5]), .QN());
   DFF_X1 \buffer_reg[9][0][1][4]  (.D(\input_filter[0][1] [4]), .CK(n_56_6), 
      .Q(\buffer[9][0][1] [4]), .QN());
   DFF_X1 \buffer_reg[9][0][1][3]  (.D(\input_filter[0][1] [3]), .CK(n_56_6), 
      .Q(\buffer[9][0][1] [3]), .QN());
   DFF_X1 \buffer_reg[9][0][1][2]  (.D(\input_filter[0][1] [2]), .CK(n_56_6), 
      .Q(\buffer[9][0][1] [2]), .QN());
   DFF_X1 \buffer_reg[9][0][1][1]  (.D(\input_filter[0][1] [1]), .CK(n_56_6), 
      .Q(\buffer[9][0][1] [1]), .QN());
   DFF_X1 \buffer_reg[9][0][1][0]  (.D(\input_filter[0][1] [0]), .CK(n_56_6), 
      .Q(\buffer[9][0][1] [0]), .QN());
   DFF_X1 \buffer_reg[10][0][1][15]  (.D(\input_filter[0][1] [15]), .CK(n_56_7), 
      .Q(\buffer[10][0][1] [15]), .QN());
   DFF_X1 \buffer_reg[10][0][1][14]  (.D(\input_filter[0][1] [14]), .CK(n_56_7), 
      .Q(\buffer[10][0][1] [14]), .QN());
   DFF_X1 \buffer_reg[10][0][1][13]  (.D(\input_filter[0][1] [13]), .CK(n_56_7), 
      .Q(\buffer[10][0][1] [13]), .QN());
   DFF_X1 \buffer_reg[10][0][1][12]  (.D(\input_filter[0][1] [12]), .CK(n_56_7), 
      .Q(\buffer[10][0][1] [12]), .QN());
   DFF_X1 \buffer_reg[10][0][1][11]  (.D(\input_filter[0][1] [11]), .CK(n_56_7), 
      .Q(\buffer[10][0][1] [11]), .QN());
   DFF_X1 \buffer_reg[10][0][1][10]  (.D(\input_filter[0][1] [10]), .CK(n_56_7), 
      .Q(\buffer[10][0][1] [10]), .QN());
   DFF_X1 \buffer_reg[10][0][1][9]  (.D(\input_filter[0][1] [9]), .CK(n_56_7), 
      .Q(\buffer[10][0][1] [9]), .QN());
   DFF_X1 \buffer_reg[10][0][1][8]  (.D(\input_filter[0][1] [8]), .CK(n_56_7), 
      .Q(\buffer[10][0][1] [8]), .QN());
   DFF_X1 \buffer_reg[10][0][1][7]  (.D(\input_filter[0][1] [7]), .CK(n_56_7), 
      .Q(\buffer[10][0][1] [7]), .QN());
   DFF_X1 \buffer_reg[10][0][1][6]  (.D(\input_filter[0][1] [6]), .CK(n_56_7), 
      .Q(\buffer[10][0][1] [6]), .QN());
   DFF_X1 \buffer_reg[10][0][1][5]  (.D(\input_filter[0][1] [5]), .CK(n_56_7), 
      .Q(\buffer[10][0][1] [5]), .QN());
   DFF_X1 \buffer_reg[10][0][1][4]  (.D(\input_filter[0][1] [4]), .CK(n_56_7), 
      .Q(\buffer[10][0][1] [4]), .QN());
   DFF_X1 \buffer_reg[10][0][1][3]  (.D(\input_filter[0][1] [3]), .CK(n_56_7), 
      .Q(\buffer[10][0][1] [3]), .QN());
   DFF_X1 \buffer_reg[10][0][1][2]  (.D(\input_filter[0][1] [2]), .CK(n_56_7), 
      .Q(\buffer[10][0][1] [2]), .QN());
   DFF_X1 \buffer_reg[10][0][1][1]  (.D(\input_filter[0][1] [1]), .CK(n_56_7), 
      .Q(\buffer[10][0][1] [1]), .QN());
   DFF_X1 \buffer_reg[10][0][1][0]  (.D(\input_filter[0][1] [0]), .CK(n_56_7), 
      .Q(\buffer[10][0][1] [0]), .QN());
   DFF_X1 \buffer_reg[11][0][1][15]  (.D(\input_filter[0][1] [15]), .CK(n_56_8), 
      .Q(\buffer[11][0][1] [15]), .QN());
   DFF_X1 \buffer_reg[11][0][1][14]  (.D(\input_filter[0][1] [14]), .CK(n_56_8), 
      .Q(\buffer[11][0][1] [14]), .QN());
   DFF_X1 \buffer_reg[11][0][1][13]  (.D(\input_filter[0][1] [13]), .CK(n_56_8), 
      .Q(\buffer[11][0][1] [13]), .QN());
   DFF_X1 \buffer_reg[11][0][1][12]  (.D(\input_filter[0][1] [12]), .CK(n_56_8), 
      .Q(\buffer[11][0][1] [12]), .QN());
   DFF_X1 \buffer_reg[11][0][1][11]  (.D(\input_filter[0][1] [11]), .CK(n_56_8), 
      .Q(\buffer[11][0][1] [11]), .QN());
   DFF_X1 \buffer_reg[11][0][1][10]  (.D(\input_filter[0][1] [10]), .CK(n_56_8), 
      .Q(\buffer[11][0][1] [10]), .QN());
   DFF_X1 \buffer_reg[11][0][1][9]  (.D(\input_filter[0][1] [9]), .CK(n_56_8), 
      .Q(\buffer[11][0][1] [9]), .QN());
   DFF_X1 \buffer_reg[11][0][1][8]  (.D(\input_filter[0][1] [8]), .CK(n_56_8), 
      .Q(\buffer[11][0][1] [8]), .QN());
   DFF_X1 \buffer_reg[11][0][1][7]  (.D(\input_filter[0][1] [7]), .CK(n_56_8), 
      .Q(\buffer[11][0][1] [7]), .QN());
   DFF_X1 \buffer_reg[11][0][1][6]  (.D(\input_filter[0][1] [6]), .CK(n_56_8), 
      .Q(\buffer[11][0][1] [6]), .QN());
   DFF_X1 \buffer_reg[11][0][1][5]  (.D(\input_filter[0][1] [5]), .CK(n_56_8), 
      .Q(\buffer[11][0][1] [5]), .QN());
   DFF_X1 \buffer_reg[11][0][1][4]  (.D(\input_filter[0][1] [4]), .CK(n_56_8), 
      .Q(\buffer[11][0][1] [4]), .QN());
   DFF_X1 \buffer_reg[11][0][1][3]  (.D(\input_filter[0][1] [3]), .CK(n_56_8), 
      .Q(\buffer[11][0][1] [3]), .QN());
   DFF_X1 \buffer_reg[11][0][1][2]  (.D(\input_filter[0][1] [2]), .CK(n_56_8), 
      .Q(\buffer[11][0][1] [2]), .QN());
   DFF_X1 \buffer_reg[11][0][1][1]  (.D(\input_filter[0][1] [1]), .CK(n_56_8), 
      .Q(\buffer[11][0][1] [1]), .QN());
   DFF_X1 \buffer_reg[11][0][1][0]  (.D(\input_filter[0][1] [0]), .CK(n_56_8), 
      .Q(\buffer[11][0][1] [0]), .QN());
   DFF_X1 \buffer_reg[12][0][1][15]  (.D(\input_filter[0][1] [15]), .CK(n_56_9), 
      .Q(\buffer[12][0][1] [15]), .QN());
   DFF_X1 \buffer_reg[12][0][1][14]  (.D(\input_filter[0][1] [14]), .CK(n_56_9), 
      .Q(\buffer[12][0][1] [14]), .QN());
   DFF_X1 \buffer_reg[12][0][1][13]  (.D(\input_filter[0][1] [13]), .CK(n_56_9), 
      .Q(\buffer[12][0][1] [13]), .QN());
   DFF_X1 \buffer_reg[12][0][1][12]  (.D(\input_filter[0][1] [12]), .CK(n_56_9), 
      .Q(\buffer[12][0][1] [12]), .QN());
   DFF_X1 \buffer_reg[12][0][1][11]  (.D(\input_filter[0][1] [11]), .CK(n_56_9), 
      .Q(\buffer[12][0][1] [11]), .QN());
   DFF_X1 \buffer_reg[12][0][1][10]  (.D(\input_filter[0][1] [10]), .CK(n_56_9), 
      .Q(\buffer[12][0][1] [10]), .QN());
   DFF_X1 \buffer_reg[12][0][1][9]  (.D(\input_filter[0][1] [9]), .CK(n_56_9), 
      .Q(\buffer[12][0][1] [9]), .QN());
   DFF_X1 \buffer_reg[12][0][1][8]  (.D(\input_filter[0][1] [8]), .CK(n_56_9), 
      .Q(\buffer[12][0][1] [8]), .QN());
   DFF_X1 \buffer_reg[12][0][1][7]  (.D(\input_filter[0][1] [7]), .CK(n_56_9), 
      .Q(\buffer[12][0][1] [7]), .QN());
   DFF_X1 \buffer_reg[12][0][1][6]  (.D(\input_filter[0][1] [6]), .CK(n_56_9), 
      .Q(\buffer[12][0][1] [6]), .QN());
   DFF_X1 \buffer_reg[12][0][1][5]  (.D(\input_filter[0][1] [5]), .CK(n_56_9), 
      .Q(\buffer[12][0][1] [5]), .QN());
   DFF_X1 \buffer_reg[12][0][1][4]  (.D(\input_filter[0][1] [4]), .CK(n_56_9), 
      .Q(\buffer[12][0][1] [4]), .QN());
   DFF_X1 \buffer_reg[12][0][1][3]  (.D(\input_filter[0][1] [3]), .CK(n_56_9), 
      .Q(\buffer[12][0][1] [3]), .QN());
   DFF_X1 \buffer_reg[12][0][1][2]  (.D(\input_filter[0][1] [2]), .CK(n_56_9), 
      .Q(\buffer[12][0][1] [2]), .QN());
   DFF_X1 \buffer_reg[12][0][1][1]  (.D(\input_filter[0][1] [1]), .CK(n_56_9), 
      .Q(\buffer[12][0][1] [1]), .QN());
   DFF_X1 \buffer_reg[12][0][1][0]  (.D(\input_filter[0][1] [0]), .CK(n_56_9), 
      .Q(\buffer[12][0][1] [0]), .QN());
   DFF_X1 \buffer_reg[13][0][1][15]  (.D(\input_filter[0][1] [15]), .CK(n_56_10), 
      .Q(\buffer[13][0][1] [15]), .QN());
   DFF_X1 \buffer_reg[13][0][1][14]  (.D(\input_filter[0][1] [14]), .CK(n_56_10), 
      .Q(\buffer[13][0][1] [14]), .QN());
   DFF_X1 \buffer_reg[13][0][1][13]  (.D(\input_filter[0][1] [13]), .CK(n_56_10), 
      .Q(\buffer[13][0][1] [13]), .QN());
   DFF_X1 \buffer_reg[13][0][1][12]  (.D(\input_filter[0][1] [12]), .CK(n_56_10), 
      .Q(\buffer[13][0][1] [12]), .QN());
   DFF_X1 \buffer_reg[13][0][1][11]  (.D(\input_filter[0][1] [11]), .CK(n_56_10), 
      .Q(\buffer[13][0][1] [11]), .QN());
   DFF_X1 \buffer_reg[13][0][1][10]  (.D(\input_filter[0][1] [10]), .CK(n_56_10), 
      .Q(\buffer[13][0][1] [10]), .QN());
   DFF_X1 \buffer_reg[13][0][1][9]  (.D(\input_filter[0][1] [9]), .CK(n_56_10), 
      .Q(\buffer[13][0][1] [9]), .QN());
   DFF_X1 \buffer_reg[13][0][1][8]  (.D(\input_filter[0][1] [8]), .CK(n_56_10), 
      .Q(\buffer[13][0][1] [8]), .QN());
   DFF_X1 \buffer_reg[13][0][1][7]  (.D(\input_filter[0][1] [7]), .CK(n_56_10), 
      .Q(\buffer[13][0][1] [7]), .QN());
   DFF_X1 \buffer_reg[13][0][1][6]  (.D(\input_filter[0][1] [6]), .CK(n_56_10), 
      .Q(\buffer[13][0][1] [6]), .QN());
   DFF_X1 \buffer_reg[13][0][1][5]  (.D(\input_filter[0][1] [5]), .CK(n_56_10), 
      .Q(\buffer[13][0][1] [5]), .QN());
   DFF_X1 \buffer_reg[13][0][1][4]  (.D(\input_filter[0][1] [4]), .CK(n_56_10), 
      .Q(\buffer[13][0][1] [4]), .QN());
   DFF_X1 \buffer_reg[13][0][1][3]  (.D(\input_filter[0][1] [3]), .CK(n_56_10), 
      .Q(\buffer[13][0][1] [3]), .QN());
   DFF_X1 \buffer_reg[13][0][1][2]  (.D(\input_filter[0][1] [2]), .CK(n_56_10), 
      .Q(\buffer[13][0][1] [2]), .QN());
   DFF_X1 \buffer_reg[13][0][1][1]  (.D(\input_filter[0][1] [1]), .CK(n_56_10), 
      .Q(\buffer[13][0][1] [1]), .QN());
   DFF_X1 \buffer_reg[13][0][1][0]  (.D(\input_filter[0][1] [0]), .CK(n_56_10), 
      .Q(\buffer[13][0][1] [0]), .QN());
   DFF_X1 \buffer_reg[14][0][1][15]  (.D(\input_filter[0][1] [15]), .CK(n_56_11), 
      .Q(\buffer[14][0][1] [15]), .QN());
   DFF_X1 \buffer_reg[14][0][1][14]  (.D(\input_filter[0][1] [14]), .CK(n_56_11), 
      .Q(\buffer[14][0][1] [14]), .QN());
   DFF_X1 \buffer_reg[14][0][1][13]  (.D(\input_filter[0][1] [13]), .CK(n_56_11), 
      .Q(\buffer[14][0][1] [13]), .QN());
   DFF_X1 \buffer_reg[14][0][1][12]  (.D(\input_filter[0][1] [12]), .CK(n_56_11), 
      .Q(\buffer[14][0][1] [12]), .QN());
   DFF_X1 \buffer_reg[14][0][1][11]  (.D(\input_filter[0][1] [11]), .CK(n_56_11), 
      .Q(\buffer[14][0][1] [11]), .QN());
   DFF_X1 \buffer_reg[14][0][1][10]  (.D(\input_filter[0][1] [10]), .CK(n_56_11), 
      .Q(\buffer[14][0][1] [10]), .QN());
   DFF_X1 \buffer_reg[14][0][1][9]  (.D(\input_filter[0][1] [9]), .CK(n_56_11), 
      .Q(\buffer[14][0][1] [9]), .QN());
   DFF_X1 \buffer_reg[14][0][1][8]  (.D(\input_filter[0][1] [8]), .CK(n_56_11), 
      .Q(\buffer[14][0][1] [8]), .QN());
   DFF_X1 \buffer_reg[14][0][1][7]  (.D(\input_filter[0][1] [7]), .CK(n_56_11), 
      .Q(\buffer[14][0][1] [7]), .QN());
   DFF_X1 \buffer_reg[14][0][1][6]  (.D(\input_filter[0][1] [6]), .CK(n_56_11), 
      .Q(\buffer[14][0][1] [6]), .QN());
   DFF_X1 \buffer_reg[14][0][1][5]  (.D(\input_filter[0][1] [5]), .CK(n_56_11), 
      .Q(\buffer[14][0][1] [5]), .QN());
   DFF_X1 \buffer_reg[14][0][1][4]  (.D(\input_filter[0][1] [4]), .CK(n_56_11), 
      .Q(\buffer[14][0][1] [4]), .QN());
   DFF_X1 \buffer_reg[14][0][1][3]  (.D(\input_filter[0][1] [3]), .CK(n_56_11), 
      .Q(\buffer[14][0][1] [3]), .QN());
   DFF_X1 \buffer_reg[14][0][1][2]  (.D(\input_filter[0][1] [2]), .CK(n_56_11), 
      .Q(\buffer[14][0][1] [2]), .QN());
   DFF_X1 \buffer_reg[14][0][1][1]  (.D(\input_filter[0][1] [1]), .CK(n_56_11), 
      .Q(\buffer[14][0][1] [1]), .QN());
   DFF_X1 \buffer_reg[14][0][1][0]  (.D(\input_filter[0][1] [0]), .CK(n_56_11), 
      .Q(\buffer[14][0][1] [0]), .QN());
   DFF_X1 \buffer_reg[15][0][1][15]  (.D(\input_filter[0][1] [15]), .CK(n_56_15), 
      .Q(\buffer[15][0][1] [15]), .QN());
   DFF_X1 \buffer_reg[15][0][1][14]  (.D(\input_filter[0][1] [14]), .CK(n_56_15), 
      .Q(\buffer[15][0][1] [14]), .QN());
   DFF_X1 \buffer_reg[15][0][1][13]  (.D(\input_filter[0][1] [13]), .CK(n_56_15), 
      .Q(\buffer[15][0][1] [13]), .QN());
   DFF_X1 \buffer_reg[15][0][1][12]  (.D(\input_filter[0][1] [12]), .CK(n_56_15), 
      .Q(\buffer[15][0][1] [12]), .QN());
   DFF_X1 \buffer_reg[15][0][1][11]  (.D(\input_filter[0][1] [11]), .CK(n_56_15), 
      .Q(\buffer[15][0][1] [11]), .QN());
   DFF_X1 \buffer_reg[15][0][1][10]  (.D(\input_filter[0][1] [10]), .CK(n_56_15), 
      .Q(\buffer[15][0][1] [10]), .QN());
   DFF_X1 \buffer_reg[15][0][1][9]  (.D(\input_filter[0][1] [9]), .CK(n_56_15), 
      .Q(\buffer[15][0][1] [9]), .QN());
   DFF_X1 \buffer_reg[15][0][1][8]  (.D(\input_filter[0][1] [8]), .CK(n_56_15), 
      .Q(\buffer[15][0][1] [8]), .QN());
   DFF_X1 \buffer_reg[15][0][1][7]  (.D(\input_filter[0][1] [7]), .CK(n_56_15), 
      .Q(\buffer[15][0][1] [7]), .QN());
   DFF_X1 \buffer_reg[15][0][1][6]  (.D(\input_filter[0][1] [6]), .CK(n_56_15), 
      .Q(\buffer[15][0][1] [6]), .QN());
   DFF_X1 \buffer_reg[15][0][1][5]  (.D(\input_filter[0][1] [5]), .CK(n_56_15), 
      .Q(\buffer[15][0][1] [5]), .QN());
   DFF_X1 \buffer_reg[15][0][1][4]  (.D(\input_filter[0][1] [4]), .CK(n_56_15), 
      .Q(\buffer[15][0][1] [4]), .QN());
   DFF_X1 \buffer_reg[15][0][1][3]  (.D(\input_filter[0][1] [3]), .CK(n_56_15), 
      .Q(\buffer[15][0][1] [3]), .QN());
   DFF_X1 \buffer_reg[15][0][1][2]  (.D(\input_filter[0][1] [2]), .CK(n_56_15), 
      .Q(\buffer[15][0][1] [2]), .QN());
   DFF_X1 \buffer_reg[15][0][1][1]  (.D(\input_filter[0][1] [1]), .CK(n_56_15), 
      .Q(\buffer[15][0][1] [1]), .QN());
   DFF_X1 \buffer_reg[15][0][1][0]  (.D(\input_filter[0][1] [0]), .CK(n_56_15), 
      .Q(\buffer[15][0][1] [0]), .QN());
   DFF_X1 \buffer_reg[6][0][2][15]  (.D(\input_filter[0][2] [15]), .CK(n_56_3), 
      .Q(\buffer[6][0][2] [15]), .QN());
   DFF_X1 \buffer_reg[6][0][2][14]  (.D(\input_filter[0][2] [14]), .CK(n_56_3), 
      .Q(\buffer[6][0][2] [14]), .QN());
   DFF_X1 \buffer_reg[6][0][2][13]  (.D(\input_filter[0][2] [13]), .CK(n_56_3), 
      .Q(\buffer[6][0][2] [13]), .QN());
   DFF_X1 \buffer_reg[6][0][2][12]  (.D(\input_filter[0][2] [12]), .CK(n_56_3), 
      .Q(\buffer[6][0][2] [12]), .QN());
   DFF_X1 \buffer_reg[6][0][2][11]  (.D(\input_filter[0][2] [11]), .CK(n_56_3), 
      .Q(\buffer[6][0][2] [11]), .QN());
   DFF_X1 \buffer_reg[6][0][2][10]  (.D(\input_filter[0][2] [10]), .CK(n_56_3), 
      .Q(\buffer[6][0][2] [10]), .QN());
   DFF_X1 \buffer_reg[6][0][2][9]  (.D(\input_filter[0][2] [9]), .CK(n_56_3), 
      .Q(\buffer[6][0][2] [9]), .QN());
   DFF_X1 \buffer_reg[6][0][2][8]  (.D(\input_filter[0][2] [8]), .CK(n_56_3), 
      .Q(\buffer[6][0][2] [8]), .QN());
   DFF_X1 \buffer_reg[6][0][2][7]  (.D(\input_filter[0][2] [7]), .CK(n_56_3), 
      .Q(\buffer[6][0][2] [7]), .QN());
   DFF_X1 \buffer_reg[6][0][2][6]  (.D(\input_filter[0][2] [6]), .CK(n_56_3), 
      .Q(\buffer[6][0][2] [6]), .QN());
   DFF_X1 \buffer_reg[6][0][2][5]  (.D(\input_filter[0][2] [5]), .CK(n_56_3), 
      .Q(\buffer[6][0][2] [5]), .QN());
   DFF_X1 \buffer_reg[6][0][2][4]  (.D(\input_filter[0][2] [4]), .CK(n_56_3), 
      .Q(\buffer[6][0][2] [4]), .QN());
   DFF_X1 \buffer_reg[6][0][2][3]  (.D(\input_filter[0][2] [3]), .CK(n_56_3), 
      .Q(\buffer[6][0][2] [3]), .QN());
   DFF_X1 \buffer_reg[6][0][2][2]  (.D(\input_filter[0][2] [2]), .CK(n_56_3), 
      .Q(\buffer[6][0][2] [2]), .QN());
   DFF_X1 \buffer_reg[6][0][2][1]  (.D(\input_filter[0][2] [1]), .CK(n_56_3), 
      .Q(\buffer[6][0][2] [1]), .QN());
   DFF_X1 \buffer_reg[6][0][2][0]  (.D(\input_filter[0][2] [0]), .CK(n_56_3), 
      .Q(\buffer[6][0][2] [0]), .QN());
   DFF_X1 \buffer_reg[15][0][2][15]  (.D(\input_filter[0][2] [15]), .CK(n_56_15), 
      .Q(\buffer[15][0][2] [15]), .QN());
   DFF_X1 \buffer_reg[15][0][2][14]  (.D(\input_filter[0][2] [14]), .CK(n_56_15), 
      .Q(\buffer[15][0][2] [14]), .QN());
   DFF_X1 \buffer_reg[15][0][2][13]  (.D(\input_filter[0][2] [13]), .CK(n_56_15), 
      .Q(\buffer[15][0][2] [13]), .QN());
   DFF_X1 \buffer_reg[15][0][2][12]  (.D(\input_filter[0][2] [12]), .CK(n_56_15), 
      .Q(\buffer[15][0][2] [12]), .QN());
   DFF_X1 \buffer_reg[15][0][2][11]  (.D(\input_filter[0][2] [11]), .CK(n_56_15), 
      .Q(\buffer[15][0][2] [11]), .QN());
   DFF_X1 \buffer_reg[15][0][2][10]  (.D(\input_filter[0][2] [10]), .CK(n_56_15), 
      .Q(\buffer[15][0][2] [10]), .QN());
   DFF_X1 \buffer_reg[15][0][2][9]  (.D(\input_filter[0][2] [9]), .CK(n_56_15), 
      .Q(\buffer[15][0][2] [9]), .QN());
   DFF_X1 \buffer_reg[15][0][2][8]  (.D(\input_filter[0][2] [8]), .CK(n_56_15), 
      .Q(\buffer[15][0][2] [8]), .QN());
   DFF_X1 \buffer_reg[15][0][2][7]  (.D(\input_filter[0][2] [7]), .CK(n_56_15), 
      .Q(\buffer[15][0][2] [7]), .QN());
   DFF_X1 \buffer_reg[15][0][2][6]  (.D(\input_filter[0][2] [6]), .CK(n_56_15), 
      .Q(\buffer[15][0][2] [6]), .QN());
   DFF_X1 \buffer_reg[15][0][2][5]  (.D(\input_filter[0][2] [5]), .CK(n_56_15), 
      .Q(\buffer[15][0][2] [5]), .QN());
   DFF_X1 \buffer_reg[15][0][2][4]  (.D(\input_filter[0][2] [4]), .CK(n_56_15), 
      .Q(\buffer[15][0][2] [4]), .QN());
   DFF_X1 \buffer_reg[15][0][2][3]  (.D(\input_filter[0][2] [3]), .CK(n_56_15), 
      .Q(\buffer[15][0][2] [3]), .QN());
   DFF_X1 \buffer_reg[15][0][2][2]  (.D(\input_filter[0][2] [2]), .CK(n_56_15), 
      .Q(\buffer[15][0][2] [2]), .QN());
   DFF_X1 \buffer_reg[15][0][2][1]  (.D(\input_filter[0][2] [1]), .CK(n_56_15), 
      .Q(\buffer[15][0][2] [1]), .QN());
   DFF_X1 \buffer_reg[15][0][2][0]  (.D(\input_filter[0][2] [0]), .CK(n_56_15), 
      .Q(\buffer[15][0][2] [0]), .QN());
   DFF_X1 \buffer_reg[1][0][3][15]  (.D(\input_filter[0][3] [15]), .CK(n_56_13), 
      .Q(\buffer[1][0][3] [15]), .QN());
   DFF_X1 \buffer_reg[1][0][3][14]  (.D(\input_filter[0][3] [14]), .CK(n_56_13), 
      .Q(\buffer[1][0][3] [14]), .QN());
   DFF_X1 \buffer_reg[1][0][3][13]  (.D(\input_filter[0][3] [13]), .CK(n_56_13), 
      .Q(\buffer[1][0][3] [13]), .QN());
   DFF_X1 \buffer_reg[1][0][3][12]  (.D(\input_filter[0][3] [12]), .CK(n_56_13), 
      .Q(\buffer[1][0][3] [12]), .QN());
   DFF_X1 \buffer_reg[1][0][3][11]  (.D(\input_filter[0][3] [11]), .CK(n_56_13), 
      .Q(\buffer[1][0][3] [11]), .QN());
   DFF_X1 \buffer_reg[1][0][3][10]  (.D(\input_filter[0][3] [10]), .CK(n_56_13), 
      .Q(\buffer[1][0][3] [10]), .QN());
   DFF_X1 \buffer_reg[1][0][3][9]  (.D(\input_filter[0][3] [9]), .CK(n_56_13), 
      .Q(\buffer[1][0][3] [9]), .QN());
   DFF_X1 \buffer_reg[1][0][3][8]  (.D(\input_filter[0][3] [8]), .CK(n_56_13), 
      .Q(\buffer[1][0][3] [8]), .QN());
   DFF_X1 \buffer_reg[1][0][3][7]  (.D(\input_filter[0][3] [7]), .CK(n_56_13), 
      .Q(\buffer[1][0][3] [7]), .QN());
   DFF_X1 \buffer_reg[1][0][3][6]  (.D(\input_filter[0][3] [6]), .CK(n_56_13), 
      .Q(\buffer[1][0][3] [6]), .QN());
   DFF_X1 \buffer_reg[1][0][3][5]  (.D(\input_filter[0][3] [5]), .CK(n_56_13), 
      .Q(\buffer[1][0][3] [5]), .QN());
   DFF_X1 \buffer_reg[1][0][3][4]  (.D(\input_filter[0][3] [4]), .CK(n_56_13), 
      .Q(\buffer[1][0][3] [4]), .QN());
   DFF_X1 \buffer_reg[1][0][3][3]  (.D(\input_filter[0][3] [3]), .CK(n_56_13), 
      .Q(\buffer[1][0][3] [3]), .QN());
   DFF_X1 \buffer_reg[1][0][3][2]  (.D(\input_filter[0][3] [2]), .CK(n_56_13), 
      .Q(\buffer[1][0][3] [2]), .QN());
   DFF_X1 \buffer_reg[1][0][3][1]  (.D(\input_filter[0][3] [1]), .CK(n_56_13), 
      .Q(\buffer[1][0][3] [1]), .QN());
   DFF_X1 \buffer_reg[1][0][3][0]  (.D(\input_filter[0][3] [0]), .CK(n_56_13), 
      .Q(\buffer[1][0][3] [0]), .QN());
   DFF_X1 \buffer_reg[2][0][3][15]  (.D(\input_filter[0][3] [15]), .CK(n_56_14), 
      .Q(\buffer[2][0][3] [15]), .QN());
   DFF_X1 \buffer_reg[2][0][3][14]  (.D(\input_filter[0][3] [14]), .CK(n_56_14), 
      .Q(\buffer[2][0][3] [14]), .QN());
   DFF_X1 \buffer_reg[2][0][3][13]  (.D(\input_filter[0][3] [13]), .CK(n_56_14), 
      .Q(\buffer[2][0][3] [13]), .QN());
   DFF_X1 \buffer_reg[2][0][3][12]  (.D(\input_filter[0][3] [12]), .CK(n_56_14), 
      .Q(\buffer[2][0][3] [12]), .QN());
   DFF_X1 \buffer_reg[2][0][3][11]  (.D(\input_filter[0][3] [11]), .CK(n_56_14), 
      .Q(\buffer[2][0][3] [11]), .QN());
   DFF_X1 \buffer_reg[2][0][3][10]  (.D(\input_filter[0][3] [10]), .CK(n_56_14), 
      .Q(\buffer[2][0][3] [10]), .QN());
   DFF_X1 \buffer_reg[2][0][3][9]  (.D(\input_filter[0][3] [9]), .CK(n_56_14), 
      .Q(\buffer[2][0][3] [9]), .QN());
   DFF_X1 \buffer_reg[2][0][3][8]  (.D(\input_filter[0][3] [8]), .CK(n_56_14), 
      .Q(\buffer[2][0][3] [8]), .QN());
   DFF_X1 \buffer_reg[2][0][3][7]  (.D(\input_filter[0][3] [7]), .CK(n_56_14), 
      .Q(\buffer[2][0][3] [7]), .QN());
   DFF_X1 \buffer_reg[2][0][3][6]  (.D(\input_filter[0][3] [6]), .CK(n_56_14), 
      .Q(\buffer[2][0][3] [6]), .QN());
   DFF_X1 \buffer_reg[2][0][3][5]  (.D(\input_filter[0][3] [5]), .CK(n_56_14), 
      .Q(\buffer[2][0][3] [5]), .QN());
   DFF_X1 \buffer_reg[2][0][3][4]  (.D(\input_filter[0][3] [4]), .CK(n_56_14), 
      .Q(\buffer[2][0][3] [4]), .QN());
   DFF_X1 \buffer_reg[2][0][3][3]  (.D(\input_filter[0][3] [3]), .CK(n_56_14), 
      .Q(\buffer[2][0][3] [3]), .QN());
   DFF_X1 \buffer_reg[2][0][3][2]  (.D(\input_filter[0][3] [2]), .CK(n_56_14), 
      .Q(\buffer[2][0][3] [2]), .QN());
   DFF_X1 \buffer_reg[2][0][3][1]  (.D(\input_filter[0][3] [1]), .CK(n_56_14), 
      .Q(\buffer[2][0][3] [1]), .QN());
   DFF_X1 \buffer_reg[2][0][3][0]  (.D(\input_filter[0][3] [0]), .CK(n_56_14), 
      .Q(\buffer[2][0][3] [0]), .QN());
   DFF_X1 \buffer_reg[3][0][3][15]  (.D(\input_filter[0][3] [15]), .CK(n_56_0), 
      .Q(\buffer[3][0][3] [15]), .QN());
   DFF_X1 \buffer_reg[3][0][3][14]  (.D(\input_filter[0][3] [14]), .CK(n_56_0), 
      .Q(\buffer[3][0][3] [14]), .QN());
   DFF_X1 \buffer_reg[3][0][3][13]  (.D(\input_filter[0][3] [13]), .CK(n_56_0), 
      .Q(\buffer[3][0][3] [13]), .QN());
   DFF_X1 \buffer_reg[3][0][3][12]  (.D(\input_filter[0][3] [12]), .CK(n_56_0), 
      .Q(\buffer[3][0][3] [12]), .QN());
   DFF_X1 \buffer_reg[3][0][3][11]  (.D(\input_filter[0][3] [11]), .CK(n_56_0), 
      .Q(\buffer[3][0][3] [11]), .QN());
   DFF_X1 \buffer_reg[3][0][3][10]  (.D(\input_filter[0][3] [10]), .CK(n_56_0), 
      .Q(\buffer[3][0][3] [10]), .QN());
   DFF_X1 \buffer_reg[3][0][3][9]  (.D(\input_filter[0][3] [9]), .CK(n_56_0), 
      .Q(\buffer[3][0][3] [9]), .QN());
   DFF_X1 \buffer_reg[3][0][3][8]  (.D(\input_filter[0][3] [8]), .CK(n_56_0), 
      .Q(\buffer[3][0][3] [8]), .QN());
   DFF_X1 \buffer_reg[3][0][3][7]  (.D(\input_filter[0][3] [7]), .CK(n_56_0), 
      .Q(\buffer[3][0][3] [7]), .QN());
   DFF_X1 \buffer_reg[3][0][3][6]  (.D(\input_filter[0][3] [6]), .CK(n_56_0), 
      .Q(\buffer[3][0][3] [6]), .QN());
   DFF_X1 \buffer_reg[3][0][3][5]  (.D(\input_filter[0][3] [5]), .CK(n_56_0), 
      .Q(\buffer[3][0][3] [5]), .QN());
   DFF_X1 \buffer_reg[3][0][3][4]  (.D(\input_filter[0][3] [4]), .CK(n_56_0), 
      .Q(\buffer[3][0][3] [4]), .QN());
   DFF_X1 \buffer_reg[3][0][3][3]  (.D(\input_filter[0][3] [3]), .CK(n_56_0), 
      .Q(\buffer[3][0][3] [3]), .QN());
   DFF_X1 \buffer_reg[3][0][3][2]  (.D(\input_filter[0][3] [2]), .CK(n_56_0), 
      .Q(\buffer[3][0][3] [2]), .QN());
   DFF_X1 \buffer_reg[3][0][3][1]  (.D(\input_filter[0][3] [1]), .CK(n_56_0), 
      .Q(\buffer[3][0][3] [1]), .QN());
   DFF_X1 \buffer_reg[3][0][3][0]  (.D(\input_filter[0][3] [0]), .CK(n_56_0), 
      .Q(\buffer[3][0][3] [0]), .QN());
   DFF_X1 \buffer_reg[10][1][4][15]  (.D(\input_filter[1][4] [15]), .CK(n_56_7), 
      .Q(\buffer[10][1][4] [15]), .QN());
   DFF_X1 \buffer_reg[10][1][4][14]  (.D(\input_filter[1][4] [14]), .CK(n_56_7), 
      .Q(\buffer[10][1][4] [14]), .QN());
   DFF_X1 \buffer_reg[10][1][4][13]  (.D(\input_filter[1][4] [13]), .CK(n_56_7), 
      .Q(\buffer[10][1][4] [13]), .QN());
   DFF_X1 \buffer_reg[10][1][4][12]  (.D(\input_filter[1][4] [12]), .CK(n_56_7), 
      .Q(\buffer[10][1][4] [12]), .QN());
   DFF_X1 \buffer_reg[10][1][4][11]  (.D(\input_filter[1][4] [11]), .CK(n_56_7), 
      .Q(\buffer[10][1][4] [11]), .QN());
   DFF_X1 \buffer_reg[10][1][4][10]  (.D(\input_filter[1][4] [10]), .CK(n_56_7), 
      .Q(\buffer[10][1][4] [10]), .QN());
   DFF_X1 \buffer_reg[10][1][4][9]  (.D(\input_filter[1][4] [9]), .CK(n_56_7), 
      .Q(\buffer[10][1][4] [9]), .QN());
   DFF_X1 \buffer_reg[10][1][4][8]  (.D(\input_filter[1][4] [8]), .CK(n_56_7), 
      .Q(\buffer[10][1][4] [8]), .QN());
   DFF_X1 \buffer_reg[10][1][4][7]  (.D(\input_filter[1][4] [7]), .CK(n_56_7), 
      .Q(\buffer[10][1][4] [7]), .QN());
   DFF_X1 \buffer_reg[10][1][4][6]  (.D(\input_filter[1][4] [6]), .CK(n_56_7), 
      .Q(\buffer[10][1][4] [6]), .QN());
   DFF_X1 \buffer_reg[10][1][4][5]  (.D(\input_filter[1][4] [5]), .CK(n_56_7), 
      .Q(\buffer[10][1][4] [5]), .QN());
   DFF_X1 \buffer_reg[10][1][4][4]  (.D(\input_filter[1][4] [4]), .CK(n_56_7), 
      .Q(\buffer[10][1][4] [4]), .QN());
   DFF_X1 \buffer_reg[10][1][4][3]  (.D(\input_filter[1][4] [3]), .CK(n_56_7), 
      .Q(\buffer[10][1][4] [3]), .QN());
   DFF_X1 \buffer_reg[10][1][4][2]  (.D(\input_filter[1][4] [2]), .CK(n_56_7), 
      .Q(\buffer[10][1][4] [2]), .QN());
   DFF_X1 \buffer_reg[10][1][4][1]  (.D(\input_filter[1][4] [1]), .CK(n_56_7), 
      .Q(\buffer[10][1][4] [1]), .QN());
   DFF_X1 \buffer_reg[10][1][4][0]  (.D(\input_filter[1][4] [0]), .CK(n_56_7), 
      .Q(\buffer[10][1][4] [0]), .QN());
   DFF_X1 \buffer_reg[9][1][4][15]  (.D(\input_filter[1][4] [15]), .CK(n_56_6), 
      .Q(\buffer[9][1][4] [15]), .QN());
   DFF_X1 \buffer_reg[9][1][4][14]  (.D(\input_filter[1][4] [14]), .CK(n_56_6), 
      .Q(\buffer[9][1][4] [14]), .QN());
   DFF_X1 \buffer_reg[9][1][4][13]  (.D(\input_filter[1][4] [13]), .CK(n_56_6), 
      .Q(\buffer[9][1][4] [13]), .QN());
   DFF_X1 \buffer_reg[9][1][4][12]  (.D(\input_filter[1][4] [12]), .CK(n_56_6), 
      .Q(\buffer[9][1][4] [12]), .QN());
   DFF_X1 \buffer_reg[9][1][4][11]  (.D(\input_filter[1][4] [11]), .CK(n_56_6), 
      .Q(\buffer[9][1][4] [11]), .QN());
   DFF_X1 \buffer_reg[9][1][4][10]  (.D(\input_filter[1][4] [10]), .CK(n_56_6), 
      .Q(\buffer[9][1][4] [10]), .QN());
   DFF_X1 \buffer_reg[9][1][4][9]  (.D(\input_filter[1][4] [9]), .CK(n_56_6), 
      .Q(\buffer[9][1][4] [9]), .QN());
   DFF_X1 \buffer_reg[9][1][4][8]  (.D(\input_filter[1][4] [8]), .CK(n_56_6), 
      .Q(\buffer[9][1][4] [8]), .QN());
   DFF_X1 \buffer_reg[9][1][4][7]  (.D(\input_filter[1][4] [7]), .CK(n_56_6), 
      .Q(\buffer[9][1][4] [7]), .QN());
   DFF_X1 \buffer_reg[9][1][4][6]  (.D(\input_filter[1][4] [6]), .CK(n_56_6), 
      .Q(\buffer[9][1][4] [6]), .QN());
   DFF_X1 \buffer_reg[9][1][4][5]  (.D(\input_filter[1][4] [5]), .CK(n_56_6), 
      .Q(\buffer[9][1][4] [5]), .QN());
   DFF_X1 \buffer_reg[9][1][4][4]  (.D(\input_filter[1][4] [4]), .CK(n_56_6), 
      .Q(\buffer[9][1][4] [4]), .QN());
   DFF_X1 \buffer_reg[9][1][4][3]  (.D(\input_filter[1][4] [3]), .CK(n_56_6), 
      .Q(\buffer[9][1][4] [3]), .QN());
   DFF_X1 \buffer_reg[9][1][4][2]  (.D(\input_filter[1][4] [2]), .CK(n_56_6), 
      .Q(\buffer[9][1][4] [2]), .QN());
   DFF_X1 \buffer_reg[9][1][4][1]  (.D(\input_filter[1][4] [1]), .CK(n_56_6), 
      .Q(\buffer[9][1][4] [1]), .QN());
   DFF_X1 \buffer_reg[9][1][4][0]  (.D(\input_filter[1][4] [0]), .CK(n_56_6), 
      .Q(\buffer[9][1][4] [0]), .QN());
   DFF_X1 \buffer_reg[8][1][4][15]  (.D(\input_filter[1][4] [15]), .CK(n_56_5), 
      .Q(\buffer[8][1][4] [15]), .QN());
   DFF_X1 \buffer_reg[8][1][4][14]  (.D(\input_filter[1][4] [14]), .CK(n_56_5), 
      .Q(\buffer[8][1][4] [14]), .QN());
   DFF_X1 \buffer_reg[8][1][4][13]  (.D(\input_filter[1][4] [13]), .CK(n_56_5), 
      .Q(\buffer[8][1][4] [13]), .QN());
   DFF_X1 \buffer_reg[8][1][4][12]  (.D(\input_filter[1][4] [12]), .CK(n_56_5), 
      .Q(\buffer[8][1][4] [12]), .QN());
   DFF_X1 \buffer_reg[8][1][4][11]  (.D(\input_filter[1][4] [11]), .CK(n_56_5), 
      .Q(\buffer[8][1][4] [11]), .QN());
   DFF_X1 \buffer_reg[8][1][4][10]  (.D(\input_filter[1][4] [10]), .CK(n_56_5), 
      .Q(\buffer[8][1][4] [10]), .QN());
   DFF_X1 \buffer_reg[8][1][4][9]  (.D(\input_filter[1][4] [9]), .CK(n_56_5), 
      .Q(\buffer[8][1][4] [9]), .QN());
   DFF_X1 \buffer_reg[8][1][4][8]  (.D(\input_filter[1][4] [8]), .CK(n_56_5), 
      .Q(\buffer[8][1][4] [8]), .QN());
   DFF_X1 \buffer_reg[8][1][4][7]  (.D(\input_filter[1][4] [7]), .CK(n_56_5), 
      .Q(\buffer[8][1][4] [7]), .QN());
   DFF_X1 \buffer_reg[8][1][4][6]  (.D(\input_filter[1][4] [6]), .CK(n_56_5), 
      .Q(\buffer[8][1][4] [6]), .QN());
   DFF_X1 \buffer_reg[8][1][4][5]  (.D(\input_filter[1][4] [5]), .CK(n_56_5), 
      .Q(\buffer[8][1][4] [5]), .QN());
   DFF_X1 \buffer_reg[8][1][4][4]  (.D(\input_filter[1][4] [4]), .CK(n_56_5), 
      .Q(\buffer[8][1][4] [4]), .QN());
   DFF_X1 \buffer_reg[8][1][4][3]  (.D(\input_filter[1][4] [3]), .CK(n_56_5), 
      .Q(\buffer[8][1][4] [3]), .QN());
   DFF_X1 \buffer_reg[8][1][4][2]  (.D(\input_filter[1][4] [2]), .CK(n_56_5), 
      .Q(\buffer[8][1][4] [2]), .QN());
   DFF_X1 \buffer_reg[8][1][4][1]  (.D(\input_filter[1][4] [1]), .CK(n_56_5), 
      .Q(\buffer[8][1][4] [1]), .QN());
   DFF_X1 \buffer_reg[8][1][4][0]  (.D(\input_filter[1][4] [0]), .CK(n_56_5), 
      .Q(\buffer[8][1][4] [0]), .QN());
   DFF_X1 \buffer_reg[7][1][4][15]  (.D(\input_filter[1][4] [15]), .CK(n_56_4), 
      .Q(\buffer[7][1][4] [15]), .QN());
   DFF_X1 \buffer_reg[7][1][4][14]  (.D(\input_filter[1][4] [14]), .CK(n_56_4), 
      .Q(\buffer[7][1][4] [14]), .QN());
   DFF_X1 \buffer_reg[7][1][4][13]  (.D(\input_filter[1][4] [13]), .CK(n_56_4), 
      .Q(\buffer[7][1][4] [13]), .QN());
   DFF_X1 \buffer_reg[7][1][4][12]  (.D(\input_filter[1][4] [12]), .CK(n_56_4), 
      .Q(\buffer[7][1][4] [12]), .QN());
   DFF_X1 \buffer_reg[7][1][4][11]  (.D(\input_filter[1][4] [11]), .CK(n_56_4), 
      .Q(\buffer[7][1][4] [11]), .QN());
   DFF_X1 \buffer_reg[7][1][4][10]  (.D(\input_filter[1][4] [10]), .CK(n_56_4), 
      .Q(\buffer[7][1][4] [10]), .QN());
   DFF_X1 \buffer_reg[7][1][4][9]  (.D(\input_filter[1][4] [9]), .CK(n_56_4), 
      .Q(\buffer[7][1][4] [9]), .QN());
   DFF_X1 \buffer_reg[7][1][4][8]  (.D(\input_filter[1][4] [8]), .CK(n_56_4), 
      .Q(\buffer[7][1][4] [8]), .QN());
   DFF_X1 \buffer_reg[7][1][4][7]  (.D(\input_filter[1][4] [7]), .CK(n_56_4), 
      .Q(\buffer[7][1][4] [7]), .QN());
   DFF_X1 \buffer_reg[7][1][4][6]  (.D(\input_filter[1][4] [6]), .CK(n_56_4), 
      .Q(\buffer[7][1][4] [6]), .QN());
   DFF_X1 \buffer_reg[7][1][4][5]  (.D(\input_filter[1][4] [5]), .CK(n_56_4), 
      .Q(\buffer[7][1][4] [5]), .QN());
   DFF_X1 \buffer_reg[7][1][4][4]  (.D(\input_filter[1][4] [4]), .CK(n_56_4), 
      .Q(\buffer[7][1][4] [4]), .QN());
   DFF_X1 \buffer_reg[7][1][4][3]  (.D(\input_filter[1][4] [3]), .CK(n_56_4), 
      .Q(\buffer[7][1][4] [3]), .QN());
   DFF_X1 \buffer_reg[7][1][4][2]  (.D(\input_filter[1][4] [2]), .CK(n_56_4), 
      .Q(\buffer[7][1][4] [2]), .QN());
   DFF_X1 \buffer_reg[7][1][4][1]  (.D(\input_filter[1][4] [1]), .CK(n_56_4), 
      .Q(\buffer[7][1][4] [1]), .QN());
   DFF_X1 \buffer_reg[7][1][4][0]  (.D(\input_filter[1][4] [0]), .CK(n_56_4), 
      .Q(\buffer[7][1][4] [0]), .QN());
   DFF_X1 \buffer_reg[6][1][4][15]  (.D(\input_filter[1][4] [15]), .CK(n_56_3), 
      .Q(\buffer[6][1][4] [15]), .QN());
   DFF_X1 \buffer_reg[6][1][4][14]  (.D(\input_filter[1][4] [14]), .CK(n_56_3), 
      .Q(\buffer[6][1][4] [14]), .QN());
   DFF_X1 \buffer_reg[6][1][4][13]  (.D(\input_filter[1][4] [13]), .CK(n_56_3), 
      .Q(\buffer[6][1][4] [13]), .QN());
   DFF_X1 \buffer_reg[6][1][4][12]  (.D(\input_filter[1][4] [12]), .CK(n_56_3), 
      .Q(\buffer[6][1][4] [12]), .QN());
   DFF_X1 \buffer_reg[6][1][4][11]  (.D(\input_filter[1][4] [11]), .CK(n_56_3), 
      .Q(\buffer[6][1][4] [11]), .QN());
   DFF_X1 \buffer_reg[6][1][4][10]  (.D(\input_filter[1][4] [10]), .CK(n_56_3), 
      .Q(\buffer[6][1][4] [10]), .QN());
   DFF_X1 \buffer_reg[6][1][4][9]  (.D(\input_filter[1][4] [9]), .CK(n_56_3), 
      .Q(\buffer[6][1][4] [9]), .QN());
   DFF_X1 \buffer_reg[6][1][4][8]  (.D(\input_filter[1][4] [8]), .CK(n_56_3), 
      .Q(\buffer[6][1][4] [8]), .QN());
   DFF_X1 \buffer_reg[6][1][4][7]  (.D(\input_filter[1][4] [7]), .CK(n_56_3), 
      .Q(\buffer[6][1][4] [7]), .QN());
   DFF_X1 \buffer_reg[6][1][4][6]  (.D(\input_filter[1][4] [6]), .CK(n_56_3), 
      .Q(\buffer[6][1][4] [6]), .QN());
   DFF_X1 \buffer_reg[6][1][4][5]  (.D(\input_filter[1][4] [5]), .CK(n_56_3), 
      .Q(\buffer[6][1][4] [5]), .QN());
   DFF_X1 \buffer_reg[6][1][4][4]  (.D(\input_filter[1][4] [4]), .CK(n_56_3), 
      .Q(\buffer[6][1][4] [4]), .QN());
   DFF_X1 \buffer_reg[6][1][4][3]  (.D(\input_filter[1][4] [3]), .CK(n_56_3), 
      .Q(\buffer[6][1][4] [3]), .QN());
   DFF_X1 \buffer_reg[6][1][4][2]  (.D(\input_filter[1][4] [2]), .CK(n_56_3), 
      .Q(\buffer[6][1][4] [2]), .QN());
   DFF_X1 \buffer_reg[6][1][4][1]  (.D(\input_filter[1][4] [1]), .CK(n_56_3), 
      .Q(\buffer[6][1][4] [1]), .QN());
   DFF_X1 \buffer_reg[6][1][4][0]  (.D(\input_filter[1][4] [0]), .CK(n_56_3), 
      .Q(\buffer[6][1][4] [0]), .QN());
   DFF_X1 \buffer_reg[5][1][4][15]  (.D(\input_filter[1][4] [15]), .CK(n_56_2), 
      .Q(\buffer[5][1][4] [15]), .QN());
   DFF_X1 \buffer_reg[5][1][4][14]  (.D(\input_filter[1][4] [14]), .CK(n_56_2), 
      .Q(\buffer[5][1][4] [14]), .QN());
   DFF_X1 \buffer_reg[5][1][4][13]  (.D(\input_filter[1][4] [13]), .CK(n_56_2), 
      .Q(\buffer[5][1][4] [13]), .QN());
   DFF_X1 \buffer_reg[5][1][4][12]  (.D(\input_filter[1][4] [12]), .CK(n_56_2), 
      .Q(\buffer[5][1][4] [12]), .QN());
   DFF_X1 \buffer_reg[5][1][4][11]  (.D(\input_filter[1][4] [11]), .CK(n_56_2), 
      .Q(\buffer[5][1][4] [11]), .QN());
   DFF_X1 \buffer_reg[5][1][4][10]  (.D(\input_filter[1][4] [10]), .CK(n_56_2), 
      .Q(\buffer[5][1][4] [10]), .QN());
   DFF_X1 \buffer_reg[5][1][4][9]  (.D(\input_filter[1][4] [9]), .CK(n_56_2), 
      .Q(\buffer[5][1][4] [9]), .QN());
   DFF_X1 \buffer_reg[5][1][4][8]  (.D(\input_filter[1][4] [8]), .CK(n_56_2), 
      .Q(\buffer[5][1][4] [8]), .QN());
   DFF_X1 \buffer_reg[5][1][4][7]  (.D(\input_filter[1][4] [7]), .CK(n_56_2), 
      .Q(\buffer[5][1][4] [7]), .QN());
   DFF_X1 \buffer_reg[5][1][4][6]  (.D(\input_filter[1][4] [6]), .CK(n_56_2), 
      .Q(\buffer[5][1][4] [6]), .QN());
   DFF_X1 \buffer_reg[5][1][4][5]  (.D(\input_filter[1][4] [5]), .CK(n_56_2), 
      .Q(\buffer[5][1][4] [5]), .QN());
   DFF_X1 \buffer_reg[5][1][4][4]  (.D(\input_filter[1][4] [4]), .CK(n_56_2), 
      .Q(\buffer[5][1][4] [4]), .QN());
   DFF_X1 \buffer_reg[5][1][4][3]  (.D(\input_filter[1][4] [3]), .CK(n_56_2), 
      .Q(\buffer[5][1][4] [3]), .QN());
   DFF_X1 \buffer_reg[5][1][4][2]  (.D(\input_filter[1][4] [2]), .CK(n_56_2), 
      .Q(\buffer[5][1][4] [2]), .QN());
   DFF_X1 \buffer_reg[5][1][4][1]  (.D(\input_filter[1][4] [1]), .CK(n_56_2), 
      .Q(\buffer[5][1][4] [1]), .QN());
   DFF_X1 \buffer_reg[5][1][4][0]  (.D(\input_filter[1][4] [0]), .CK(n_56_2), 
      .Q(\buffer[5][1][4] [0]), .QN());
   DFF_X1 \buffer_reg[4][1][4][15]  (.D(\input_filter[1][4] [15]), .CK(n_56_1), 
      .Q(\buffer[4][1][4] [15]), .QN());
   DFF_X1 \buffer_reg[4][1][4][14]  (.D(\input_filter[1][4] [14]), .CK(n_56_1), 
      .Q(\buffer[4][1][4] [14]), .QN());
   DFF_X1 \buffer_reg[4][1][4][13]  (.D(\input_filter[1][4] [13]), .CK(n_56_1), 
      .Q(\buffer[4][1][4] [13]), .QN());
   DFF_X1 \buffer_reg[4][1][4][12]  (.D(\input_filter[1][4] [12]), .CK(n_56_1), 
      .Q(\buffer[4][1][4] [12]), .QN());
   DFF_X1 \buffer_reg[4][1][4][11]  (.D(\input_filter[1][4] [11]), .CK(n_56_1), 
      .Q(\buffer[4][1][4] [11]), .QN());
   DFF_X1 \buffer_reg[4][1][4][10]  (.D(\input_filter[1][4] [10]), .CK(n_56_1), 
      .Q(\buffer[4][1][4] [10]), .QN());
   DFF_X1 \buffer_reg[4][1][4][9]  (.D(\input_filter[1][4] [9]), .CK(n_56_1), 
      .Q(\buffer[4][1][4] [9]), .QN());
   DFF_X1 \buffer_reg[4][1][4][8]  (.D(\input_filter[1][4] [8]), .CK(n_56_1), 
      .Q(\buffer[4][1][4] [8]), .QN());
   DFF_X1 \buffer_reg[4][1][4][7]  (.D(\input_filter[1][4] [7]), .CK(n_56_1), 
      .Q(\buffer[4][1][4] [7]), .QN());
   DFF_X1 \buffer_reg[4][1][4][6]  (.D(\input_filter[1][4] [6]), .CK(n_56_1), 
      .Q(\buffer[4][1][4] [6]), .QN());
   DFF_X1 \buffer_reg[4][1][4][5]  (.D(\input_filter[1][4] [5]), .CK(n_56_1), 
      .Q(\buffer[4][1][4] [5]), .QN());
   DFF_X1 \buffer_reg[4][1][4][4]  (.D(\input_filter[1][4] [4]), .CK(n_56_1), 
      .Q(\buffer[4][1][4] [4]), .QN());
   DFF_X1 \buffer_reg[4][1][4][3]  (.D(\input_filter[1][4] [3]), .CK(n_56_1), 
      .Q(\buffer[4][1][4] [3]), .QN());
   DFF_X1 \buffer_reg[4][1][4][2]  (.D(\input_filter[1][4] [2]), .CK(n_56_1), 
      .Q(\buffer[4][1][4] [2]), .QN());
   DFF_X1 \buffer_reg[4][1][4][1]  (.D(\input_filter[1][4] [1]), .CK(n_56_1), 
      .Q(\buffer[4][1][4] [1]), .QN());
   DFF_X1 \buffer_reg[4][1][4][0]  (.D(\input_filter[1][4] [0]), .CK(n_56_1), 
      .Q(\buffer[4][1][4] [0]), .QN());
   DFF_X1 \buffer_reg[3][1][4][15]  (.D(\input_filter[1][4] [15]), .CK(n_56_0), 
      .Q(\buffer[3][1][4] [15]), .QN());
   DFF_X1 \buffer_reg[3][1][4][14]  (.D(\input_filter[1][4] [14]), .CK(n_56_0), 
      .Q(\buffer[3][1][4] [14]), .QN());
   DFF_X1 \buffer_reg[3][1][4][13]  (.D(\input_filter[1][4] [13]), .CK(n_56_0), 
      .Q(\buffer[3][1][4] [13]), .QN());
   DFF_X1 \buffer_reg[3][1][4][12]  (.D(\input_filter[1][4] [12]), .CK(n_56_0), 
      .Q(\buffer[3][1][4] [12]), .QN());
   DFF_X1 \buffer_reg[3][1][4][11]  (.D(\input_filter[1][4] [11]), .CK(n_56_0), 
      .Q(\buffer[3][1][4] [11]), .QN());
   DFF_X1 \buffer_reg[3][1][4][10]  (.D(\input_filter[1][4] [10]), .CK(n_56_0), 
      .Q(\buffer[3][1][4] [10]), .QN());
   DFF_X1 \buffer_reg[3][1][4][9]  (.D(\input_filter[1][4] [9]), .CK(n_56_0), 
      .Q(\buffer[3][1][4] [9]), .QN());
   DFF_X1 \buffer_reg[3][1][4][8]  (.D(\input_filter[1][4] [8]), .CK(n_56_0), 
      .Q(\buffer[3][1][4] [8]), .QN());
   DFF_X1 \buffer_reg[3][1][4][7]  (.D(\input_filter[1][4] [7]), .CK(n_56_0), 
      .Q(\buffer[3][1][4] [7]), .QN());
   DFF_X1 \buffer_reg[3][1][4][6]  (.D(\input_filter[1][4] [6]), .CK(n_56_0), 
      .Q(\buffer[3][1][4] [6]), .QN());
   DFF_X1 \buffer_reg[3][1][4][5]  (.D(\input_filter[1][4] [5]), .CK(n_56_0), 
      .Q(\buffer[3][1][4] [5]), .QN());
   DFF_X1 \buffer_reg[3][1][4][4]  (.D(\input_filter[1][4] [4]), .CK(n_56_0), 
      .Q(\buffer[3][1][4] [4]), .QN());
   DFF_X1 \buffer_reg[3][1][4][3]  (.D(\input_filter[1][4] [3]), .CK(n_56_0), 
      .Q(\buffer[3][1][4] [3]), .QN());
   DFF_X1 \buffer_reg[3][1][4][2]  (.D(\input_filter[1][4] [2]), .CK(n_56_0), 
      .Q(\buffer[3][1][4] [2]), .QN());
   DFF_X1 \buffer_reg[3][1][4][1]  (.D(\input_filter[1][4] [1]), .CK(n_56_0), 
      .Q(\buffer[3][1][4] [1]), .QN());
   DFF_X1 \buffer_reg[3][1][4][0]  (.D(\input_filter[1][4] [0]), .CK(n_56_0), 
      .Q(\buffer[3][1][4] [0]), .QN());
   DFF_X1 \buffer_reg[2][1][4][15]  (.D(\input_filter[1][4] [15]), .CK(n_56_14), 
      .Q(\buffer[2][1][4] [15]), .QN());
   DFF_X1 \buffer_reg[2][1][4][14]  (.D(\input_filter[1][4] [14]), .CK(n_56_14), 
      .Q(\buffer[2][1][4] [14]), .QN());
   DFF_X1 \buffer_reg[2][1][4][13]  (.D(\input_filter[1][4] [13]), .CK(n_56_14), 
      .Q(\buffer[2][1][4] [13]), .QN());
   DFF_X1 \buffer_reg[2][1][4][12]  (.D(\input_filter[1][4] [12]), .CK(n_56_14), 
      .Q(\buffer[2][1][4] [12]), .QN());
   DFF_X1 \buffer_reg[2][1][4][11]  (.D(\input_filter[1][4] [11]), .CK(n_56_14), 
      .Q(\buffer[2][1][4] [11]), .QN());
   DFF_X1 \buffer_reg[2][1][4][10]  (.D(\input_filter[1][4] [10]), .CK(n_56_14), 
      .Q(\buffer[2][1][4] [10]), .QN());
   DFF_X1 \buffer_reg[2][1][4][9]  (.D(\input_filter[1][4] [9]), .CK(n_56_14), 
      .Q(\buffer[2][1][4] [9]), .QN());
   DFF_X1 \buffer_reg[2][1][4][8]  (.D(\input_filter[1][4] [8]), .CK(n_56_14), 
      .Q(\buffer[2][1][4] [8]), .QN());
   DFF_X1 \buffer_reg[2][1][4][7]  (.D(\input_filter[1][4] [7]), .CK(n_56_14), 
      .Q(\buffer[2][1][4] [7]), .QN());
   DFF_X1 \buffer_reg[2][1][4][6]  (.D(\input_filter[1][4] [6]), .CK(n_56_14), 
      .Q(\buffer[2][1][4] [6]), .QN());
   DFF_X1 \buffer_reg[2][1][4][5]  (.D(\input_filter[1][4] [5]), .CK(n_56_14), 
      .Q(\buffer[2][1][4] [5]), .QN());
   DFF_X1 \buffer_reg[2][1][4][4]  (.D(\input_filter[1][4] [4]), .CK(n_56_14), 
      .Q(\buffer[2][1][4] [4]), .QN());
   DFF_X1 \buffer_reg[2][1][4][3]  (.D(\input_filter[1][4] [3]), .CK(n_56_14), 
      .Q(\buffer[2][1][4] [3]), .QN());
   DFF_X1 \buffer_reg[2][1][4][2]  (.D(\input_filter[1][4] [2]), .CK(n_56_14), 
      .Q(\buffer[2][1][4] [2]), .QN());
   DFF_X1 \buffer_reg[2][1][4][1]  (.D(\input_filter[1][4] [1]), .CK(n_56_14), 
      .Q(\buffer[2][1][4] [1]), .QN());
   DFF_X1 \buffer_reg[2][1][4][0]  (.D(\input_filter[1][4] [0]), .CK(n_56_14), 
      .Q(\buffer[2][1][4] [0]), .QN());
   DFF_X1 \buffer_reg[1][1][4][15]  (.D(\input_filter[1][4] [15]), .CK(n_56_13), 
      .Q(\buffer[1][1][4] [15]), .QN());
   DFF_X1 \buffer_reg[1][1][4][14]  (.D(\input_filter[1][4] [14]), .CK(n_56_13), 
      .Q(\buffer[1][1][4] [14]), .QN());
   DFF_X1 \buffer_reg[1][1][4][13]  (.D(\input_filter[1][4] [13]), .CK(n_56_13), 
      .Q(\buffer[1][1][4] [13]), .QN());
   DFF_X1 \buffer_reg[1][1][4][12]  (.D(\input_filter[1][4] [12]), .CK(n_56_13), 
      .Q(\buffer[1][1][4] [12]), .QN());
   DFF_X1 \buffer_reg[1][1][4][11]  (.D(\input_filter[1][4] [11]), .CK(n_56_13), 
      .Q(\buffer[1][1][4] [11]), .QN());
   DFF_X1 \buffer_reg[1][1][4][10]  (.D(\input_filter[1][4] [10]), .CK(n_56_13), 
      .Q(\buffer[1][1][4] [10]), .QN());
   DFF_X1 \buffer_reg[1][1][4][9]  (.D(\input_filter[1][4] [9]), .CK(n_56_13), 
      .Q(\buffer[1][1][4] [9]), .QN());
   DFF_X1 \buffer_reg[1][1][4][8]  (.D(\input_filter[1][4] [8]), .CK(n_56_13), 
      .Q(\buffer[1][1][4] [8]), .QN());
   DFF_X1 \buffer_reg[1][1][4][7]  (.D(\input_filter[1][4] [7]), .CK(n_56_13), 
      .Q(\buffer[1][1][4] [7]), .QN());
   DFF_X1 \buffer_reg[1][1][4][6]  (.D(\input_filter[1][4] [6]), .CK(n_56_13), 
      .Q(\buffer[1][1][4] [6]), .QN());
   DFF_X1 \buffer_reg[1][1][4][5]  (.D(\input_filter[1][4] [5]), .CK(n_56_13), 
      .Q(\buffer[1][1][4] [5]), .QN());
   DFF_X1 \buffer_reg[1][1][4][4]  (.D(\input_filter[1][4] [4]), .CK(n_56_13), 
      .Q(\buffer[1][1][4] [4]), .QN());
   DFF_X1 \buffer_reg[1][1][4][3]  (.D(\input_filter[1][4] [3]), .CK(n_56_13), 
      .Q(\buffer[1][1][4] [3]), .QN());
   DFF_X1 \buffer_reg[1][1][4][2]  (.D(\input_filter[1][4] [2]), .CK(n_56_13), 
      .Q(\buffer[1][1][4] [2]), .QN());
   DFF_X1 \buffer_reg[1][1][4][1]  (.D(\input_filter[1][4] [1]), .CK(n_56_13), 
      .Q(\buffer[1][1][4] [1]), .QN());
   DFF_X1 \buffer_reg[1][1][4][0]  (.D(\input_filter[1][4] [0]), .CK(n_56_13), 
      .Q(\buffer[1][1][4] [0]), .QN());
   DFF_X1 \buffer_reg[4][0][3][15]  (.D(\input_filter[0][3] [15]), .CK(n_56_1), 
      .Q(\buffer[4][0][3] [15]), .QN());
   DFF_X1 \buffer_reg[4][0][3][14]  (.D(\input_filter[0][3] [14]), .CK(n_56_1), 
      .Q(\buffer[4][0][3] [14]), .QN());
   DFF_X1 \buffer_reg[4][0][3][13]  (.D(\input_filter[0][3] [13]), .CK(n_56_1), 
      .Q(\buffer[4][0][3] [13]), .QN());
   DFF_X1 \buffer_reg[4][0][3][12]  (.D(\input_filter[0][3] [12]), .CK(n_56_1), 
      .Q(\buffer[4][0][3] [12]), .QN());
   DFF_X1 \buffer_reg[4][0][3][11]  (.D(\input_filter[0][3] [11]), .CK(n_56_1), 
      .Q(\buffer[4][0][3] [11]), .QN());
   DFF_X1 \buffer_reg[4][0][3][10]  (.D(\input_filter[0][3] [10]), .CK(n_56_1), 
      .Q(\buffer[4][0][3] [10]), .QN());
   DFF_X1 \buffer_reg[4][0][3][9]  (.D(\input_filter[0][3] [9]), .CK(n_56_1), 
      .Q(\buffer[4][0][3] [9]), .QN());
   DFF_X1 \buffer_reg[4][0][3][8]  (.D(\input_filter[0][3] [8]), .CK(n_56_1), 
      .Q(\buffer[4][0][3] [8]), .QN());
   DFF_X1 \buffer_reg[4][0][3][7]  (.D(\input_filter[0][3] [7]), .CK(n_56_1), 
      .Q(\buffer[4][0][3] [7]), .QN());
   DFF_X1 \buffer_reg[4][0][3][6]  (.D(\input_filter[0][3] [6]), .CK(n_56_1), 
      .Q(\buffer[4][0][3] [6]), .QN());
   DFF_X1 \buffer_reg[4][0][3][5]  (.D(\input_filter[0][3] [5]), .CK(n_56_1), 
      .Q(\buffer[4][0][3] [5]), .QN());
   DFF_X1 \buffer_reg[4][0][3][4]  (.D(\input_filter[0][3] [4]), .CK(n_56_1), 
      .Q(\buffer[4][0][3] [4]), .QN());
   DFF_X1 \buffer_reg[4][0][3][3]  (.D(\input_filter[0][3] [3]), .CK(n_56_1), 
      .Q(\buffer[4][0][3] [3]), .QN());
   DFF_X1 \buffer_reg[4][0][3][2]  (.D(\input_filter[0][3] [2]), .CK(n_56_1), 
      .Q(\buffer[4][0][3] [2]), .QN());
   DFF_X1 \buffer_reg[4][0][3][1]  (.D(\input_filter[0][3] [1]), .CK(n_56_1), 
      .Q(\buffer[4][0][3] [1]), .QN());
   DFF_X1 \buffer_reg[4][0][3][0]  (.D(\input_filter[0][3] [0]), .CK(n_56_1), 
      .Q(\buffer[4][0][3] [0]), .QN());
   DFF_X1 \buffer_reg[5][0][3][15]  (.D(\input_filter[0][3] [15]), .CK(n_56_2), 
      .Q(\buffer[5][0][3] [15]), .QN());
   DFF_X1 \buffer_reg[5][0][3][14]  (.D(\input_filter[0][3] [14]), .CK(n_56_2), 
      .Q(\buffer[5][0][3] [14]), .QN());
   DFF_X1 \buffer_reg[5][0][3][13]  (.D(\input_filter[0][3] [13]), .CK(n_56_2), 
      .Q(\buffer[5][0][3] [13]), .QN());
   DFF_X1 \buffer_reg[5][0][3][12]  (.D(\input_filter[0][3] [12]), .CK(n_56_2), 
      .Q(\buffer[5][0][3] [12]), .QN());
   DFF_X1 \buffer_reg[5][0][3][11]  (.D(\input_filter[0][3] [11]), .CK(n_56_2), 
      .Q(\buffer[5][0][3] [11]), .QN());
   DFF_X1 \buffer_reg[5][0][3][10]  (.D(\input_filter[0][3] [10]), .CK(n_56_2), 
      .Q(\buffer[5][0][3] [10]), .QN());
   DFF_X1 \buffer_reg[5][0][3][9]  (.D(\input_filter[0][3] [9]), .CK(n_56_2), 
      .Q(\buffer[5][0][3] [9]), .QN());
   DFF_X1 \buffer_reg[5][0][3][8]  (.D(\input_filter[0][3] [8]), .CK(n_56_2), 
      .Q(\buffer[5][0][3] [8]), .QN());
   DFF_X1 \buffer_reg[5][0][3][7]  (.D(\input_filter[0][3] [7]), .CK(n_56_2), 
      .Q(\buffer[5][0][3] [7]), .QN());
   DFF_X1 \buffer_reg[5][0][3][6]  (.D(\input_filter[0][3] [6]), .CK(n_56_2), 
      .Q(\buffer[5][0][3] [6]), .QN());
   DFF_X1 \buffer_reg[5][0][3][5]  (.D(\input_filter[0][3] [5]), .CK(n_56_2), 
      .Q(\buffer[5][0][3] [5]), .QN());
   DFF_X1 \buffer_reg[5][0][3][4]  (.D(\input_filter[0][3] [4]), .CK(n_56_2), 
      .Q(\buffer[5][0][3] [4]), .QN());
   DFF_X1 \buffer_reg[5][0][3][3]  (.D(\input_filter[0][3] [3]), .CK(n_56_2), 
      .Q(\buffer[5][0][3] [3]), .QN());
   DFF_X1 \buffer_reg[5][0][3][2]  (.D(\input_filter[0][3] [2]), .CK(n_56_2), 
      .Q(\buffer[5][0][3] [2]), .QN());
   DFF_X1 \buffer_reg[5][0][3][1]  (.D(\input_filter[0][3] [1]), .CK(n_56_2), 
      .Q(\buffer[5][0][3] [1]), .QN());
   DFF_X1 \buffer_reg[5][0][3][0]  (.D(\input_filter[0][3] [0]), .CK(n_56_2), 
      .Q(\buffer[5][0][3] [0]), .QN());
   DFF_X1 \buffer_reg[6][0][3][15]  (.D(\input_filter[0][3] [15]), .CK(n_56_3), 
      .Q(\buffer[6][0][3] [15]), .QN());
   DFF_X1 \buffer_reg[6][0][3][14]  (.D(\input_filter[0][3] [14]), .CK(n_56_3), 
      .Q(\buffer[6][0][3] [14]), .QN());
   DFF_X1 \buffer_reg[6][0][3][13]  (.D(\input_filter[0][3] [13]), .CK(n_56_3), 
      .Q(\buffer[6][0][3] [13]), .QN());
   DFF_X1 \buffer_reg[6][0][3][12]  (.D(\input_filter[0][3] [12]), .CK(n_56_3), 
      .Q(\buffer[6][0][3] [12]), .QN());
   DFF_X1 \buffer_reg[6][0][3][11]  (.D(\input_filter[0][3] [11]), .CK(n_56_3), 
      .Q(\buffer[6][0][3] [11]), .QN());
   DFF_X1 \buffer_reg[6][0][3][10]  (.D(\input_filter[0][3] [10]), .CK(n_56_3), 
      .Q(\buffer[6][0][3] [10]), .QN());
   DFF_X1 \buffer_reg[6][0][3][9]  (.D(\input_filter[0][3] [9]), .CK(n_56_3), 
      .Q(\buffer[6][0][3] [9]), .QN());
   DFF_X1 \buffer_reg[6][0][3][8]  (.D(\input_filter[0][3] [8]), .CK(n_56_3), 
      .Q(\buffer[6][0][3] [8]), .QN());
   DFF_X1 \buffer_reg[6][0][3][7]  (.D(\input_filter[0][3] [7]), .CK(n_56_3), 
      .Q(\buffer[6][0][3] [7]), .QN());
   DFF_X1 \buffer_reg[6][0][3][6]  (.D(\input_filter[0][3] [6]), .CK(n_56_3), 
      .Q(\buffer[6][0][3] [6]), .QN());
   DFF_X1 \buffer_reg[6][0][3][5]  (.D(\input_filter[0][3] [5]), .CK(n_56_3), 
      .Q(\buffer[6][0][3] [5]), .QN());
   DFF_X1 \buffer_reg[6][0][3][4]  (.D(\input_filter[0][3] [4]), .CK(n_56_3), 
      .Q(\buffer[6][0][3] [4]), .QN());
   DFF_X1 \buffer_reg[6][0][3][3]  (.D(\input_filter[0][3] [3]), .CK(n_56_3), 
      .Q(\buffer[6][0][3] [3]), .QN());
   DFF_X1 \buffer_reg[6][0][3][2]  (.D(\input_filter[0][3] [2]), .CK(n_56_3), 
      .Q(\buffer[6][0][3] [2]), .QN());
   DFF_X1 \buffer_reg[6][0][3][1]  (.D(\input_filter[0][3] [1]), .CK(n_56_3), 
      .Q(\buffer[6][0][3] [1]), .QN());
   DFF_X1 \buffer_reg[6][0][3][0]  (.D(\input_filter[0][3] [0]), .CK(n_56_3), 
      .Q(\buffer[6][0][3] [0]), .QN());
   DFF_X1 \buffer_reg[7][0][3][15]  (.D(\input_filter[0][3] [15]), .CK(n_56_4), 
      .Q(\buffer[7][0][3] [15]), .QN());
   DFF_X1 \buffer_reg[7][0][3][14]  (.D(\input_filter[0][3] [14]), .CK(n_56_4), 
      .Q(\buffer[7][0][3] [14]), .QN());
   DFF_X1 \buffer_reg[7][0][3][13]  (.D(\input_filter[0][3] [13]), .CK(n_56_4), 
      .Q(\buffer[7][0][3] [13]), .QN());
   DFF_X1 \buffer_reg[7][0][3][12]  (.D(\input_filter[0][3] [12]), .CK(n_56_4), 
      .Q(\buffer[7][0][3] [12]), .QN());
   DFF_X1 \buffer_reg[7][0][3][11]  (.D(\input_filter[0][3] [11]), .CK(n_56_4), 
      .Q(\buffer[7][0][3] [11]), .QN());
   DFF_X1 \buffer_reg[7][0][3][10]  (.D(\input_filter[0][3] [10]), .CK(n_56_4), 
      .Q(\buffer[7][0][3] [10]), .QN());
   DFF_X1 \buffer_reg[7][0][3][9]  (.D(\input_filter[0][3] [9]), .CK(n_56_4), 
      .Q(\buffer[7][0][3] [9]), .QN());
   DFF_X1 \buffer_reg[7][0][3][8]  (.D(\input_filter[0][3] [8]), .CK(n_56_4), 
      .Q(\buffer[7][0][3] [8]), .QN());
   DFF_X1 \buffer_reg[7][0][3][7]  (.D(\input_filter[0][3] [7]), .CK(n_56_4), 
      .Q(\buffer[7][0][3] [7]), .QN());
   DFF_X1 \buffer_reg[7][0][3][6]  (.D(\input_filter[0][3] [6]), .CK(n_56_4), 
      .Q(\buffer[7][0][3] [6]), .QN());
   DFF_X1 \buffer_reg[7][0][3][5]  (.D(\input_filter[0][3] [5]), .CK(n_56_4), 
      .Q(\buffer[7][0][3] [5]), .QN());
   DFF_X1 \buffer_reg[7][0][3][4]  (.D(\input_filter[0][3] [4]), .CK(n_56_4), 
      .Q(\buffer[7][0][3] [4]), .QN());
   DFF_X1 \buffer_reg[7][0][3][3]  (.D(\input_filter[0][3] [3]), .CK(n_56_4), 
      .Q(\buffer[7][0][3] [3]), .QN());
   DFF_X1 \buffer_reg[7][0][3][2]  (.D(\input_filter[0][3] [2]), .CK(n_56_4), 
      .Q(\buffer[7][0][3] [2]), .QN());
   DFF_X1 \buffer_reg[7][0][3][1]  (.D(\input_filter[0][3] [1]), .CK(n_56_4), 
      .Q(\buffer[7][0][3] [1]), .QN());
   DFF_X1 \buffer_reg[7][0][3][0]  (.D(\input_filter[0][3] [0]), .CK(n_56_4), 
      .Q(\buffer[7][0][3] [0]), .QN());
   DFF_X1 \buffer_reg[8][0][3][15]  (.D(\input_filter[0][3] [15]), .CK(n_56_5), 
      .Q(\buffer[8][0][3] [15]), .QN());
   DFF_X1 \buffer_reg[8][0][3][14]  (.D(\input_filter[0][3] [14]), .CK(n_56_5), 
      .Q(\buffer[8][0][3] [14]), .QN());
   DFF_X1 \buffer_reg[8][0][3][13]  (.D(\input_filter[0][3] [13]), .CK(n_56_5), 
      .Q(\buffer[8][0][3] [13]), .QN());
   DFF_X1 \buffer_reg[8][0][3][12]  (.D(\input_filter[0][3] [12]), .CK(n_56_5), 
      .Q(\buffer[8][0][3] [12]), .QN());
   DFF_X1 \buffer_reg[8][0][3][11]  (.D(\input_filter[0][3] [11]), .CK(n_56_5), 
      .Q(\buffer[8][0][3] [11]), .QN());
   DFF_X1 \buffer_reg[8][0][3][10]  (.D(\input_filter[0][3] [10]), .CK(n_56_5), 
      .Q(\buffer[8][0][3] [10]), .QN());
   DFF_X1 \buffer_reg[8][0][3][9]  (.D(\input_filter[0][3] [9]), .CK(n_56_5), 
      .Q(\buffer[8][0][3] [9]), .QN());
   DFF_X1 \buffer_reg[8][0][3][8]  (.D(\input_filter[0][3] [8]), .CK(n_56_5), 
      .Q(\buffer[8][0][3] [8]), .QN());
   DFF_X1 \buffer_reg[8][0][3][7]  (.D(\input_filter[0][3] [7]), .CK(n_56_5), 
      .Q(\buffer[8][0][3] [7]), .QN());
   DFF_X1 \buffer_reg[8][0][3][6]  (.D(\input_filter[0][3] [6]), .CK(n_56_5), 
      .Q(\buffer[8][0][3] [6]), .QN());
   DFF_X1 \buffer_reg[8][0][3][5]  (.D(\input_filter[0][3] [5]), .CK(n_56_5), 
      .Q(\buffer[8][0][3] [5]), .QN());
   DFF_X1 \buffer_reg[8][0][3][4]  (.D(\input_filter[0][3] [4]), .CK(n_56_5), 
      .Q(\buffer[8][0][3] [4]), .QN());
   DFF_X1 \buffer_reg[8][0][3][3]  (.D(\input_filter[0][3] [3]), .CK(n_56_5), 
      .Q(\buffer[8][0][3] [3]), .QN());
   DFF_X1 \buffer_reg[8][0][3][2]  (.D(\input_filter[0][3] [2]), .CK(n_56_5), 
      .Q(\buffer[8][0][3] [2]), .QN());
   DFF_X1 \buffer_reg[8][0][3][1]  (.D(\input_filter[0][3] [1]), .CK(n_56_5), 
      .Q(\buffer[8][0][3] [1]), .QN());
   DFF_X1 \buffer_reg[8][0][3][0]  (.D(\input_filter[0][3] [0]), .CK(n_56_5), 
      .Q(\buffer[8][0][3] [0]), .QN());
   DFF_X1 \buffer_reg[9][0][3][15]  (.D(\input_filter[0][3] [15]), .CK(n_56_6), 
      .Q(\buffer[9][0][3] [15]), .QN());
   DFF_X1 \buffer_reg[9][0][3][14]  (.D(\input_filter[0][3] [14]), .CK(n_56_6), 
      .Q(\buffer[9][0][3] [14]), .QN());
   DFF_X1 \buffer_reg[9][0][3][13]  (.D(\input_filter[0][3] [13]), .CK(n_56_6), 
      .Q(\buffer[9][0][3] [13]), .QN());
   DFF_X1 \buffer_reg[9][0][3][12]  (.D(\input_filter[0][3] [12]), .CK(n_56_6), 
      .Q(\buffer[9][0][3] [12]), .QN());
   DFF_X1 \buffer_reg[9][0][3][11]  (.D(\input_filter[0][3] [11]), .CK(n_56_6), 
      .Q(\buffer[9][0][3] [11]), .QN());
   DFF_X1 \buffer_reg[9][0][3][10]  (.D(\input_filter[0][3] [10]), .CK(n_56_6), 
      .Q(\buffer[9][0][3] [10]), .QN());
   DFF_X1 \buffer_reg[9][0][3][9]  (.D(\input_filter[0][3] [9]), .CK(n_56_6), 
      .Q(\buffer[9][0][3] [9]), .QN());
   DFF_X1 \buffer_reg[9][0][3][8]  (.D(\input_filter[0][3] [8]), .CK(n_56_6), 
      .Q(\buffer[9][0][3] [8]), .QN());
   DFF_X1 \buffer_reg[9][0][3][7]  (.D(\input_filter[0][3] [7]), .CK(n_56_6), 
      .Q(\buffer[9][0][3] [7]), .QN());
   DFF_X1 \buffer_reg[9][0][3][6]  (.D(\input_filter[0][3] [6]), .CK(n_56_6), 
      .Q(\buffer[9][0][3] [6]), .QN());
   DFF_X1 \buffer_reg[9][0][3][5]  (.D(\input_filter[0][3] [5]), .CK(n_56_6), 
      .Q(\buffer[9][0][3] [5]), .QN());
   DFF_X1 \buffer_reg[9][0][3][4]  (.D(\input_filter[0][3] [4]), .CK(n_56_6), 
      .Q(\buffer[9][0][3] [4]), .QN());
   DFF_X1 \buffer_reg[9][0][3][3]  (.D(\input_filter[0][3] [3]), .CK(n_56_6), 
      .Q(\buffer[9][0][3] [3]), .QN());
   DFF_X1 \buffer_reg[9][0][3][2]  (.D(\input_filter[0][3] [2]), .CK(n_56_6), 
      .Q(\buffer[9][0][3] [2]), .QN());
   DFF_X1 \buffer_reg[9][0][3][1]  (.D(\input_filter[0][3] [1]), .CK(n_56_6), 
      .Q(\buffer[9][0][3] [1]), .QN());
   DFF_X1 \buffer_reg[9][0][3][0]  (.D(\input_filter[0][3] [0]), .CK(n_56_6), 
      .Q(\buffer[9][0][3] [0]), .QN());
   DFF_X1 \buffer_reg[10][0][3][15]  (.D(\input_filter[0][3] [15]), .CK(n_56_7), 
      .Q(\buffer[10][0][3] [15]), .QN());
   DFF_X1 \buffer_reg[10][0][3][14]  (.D(\input_filter[0][3] [14]), .CK(n_56_7), 
      .Q(\buffer[10][0][3] [14]), .QN());
   DFF_X1 \buffer_reg[10][0][3][13]  (.D(\input_filter[0][3] [13]), .CK(n_56_7), 
      .Q(\buffer[10][0][3] [13]), .QN());
   DFF_X1 \buffer_reg[10][0][3][12]  (.D(\input_filter[0][3] [12]), .CK(n_56_7), 
      .Q(\buffer[10][0][3] [12]), .QN());
   DFF_X1 \buffer_reg[10][0][3][11]  (.D(\input_filter[0][3] [11]), .CK(n_56_7), 
      .Q(\buffer[10][0][3] [11]), .QN());
   DFF_X1 \buffer_reg[10][0][3][10]  (.D(\input_filter[0][3] [10]), .CK(n_56_7), 
      .Q(\buffer[10][0][3] [10]), .QN());
   DFF_X1 \buffer_reg[10][0][3][9]  (.D(\input_filter[0][3] [9]), .CK(n_56_7), 
      .Q(\buffer[10][0][3] [9]), .QN());
   DFF_X1 \buffer_reg[10][0][3][8]  (.D(\input_filter[0][3] [8]), .CK(n_56_7), 
      .Q(\buffer[10][0][3] [8]), .QN());
   DFF_X1 \buffer_reg[10][0][3][7]  (.D(\input_filter[0][3] [7]), .CK(n_56_7), 
      .Q(\buffer[10][0][3] [7]), .QN());
   DFF_X1 \buffer_reg[10][0][3][6]  (.D(\input_filter[0][3] [6]), .CK(n_56_7), 
      .Q(\buffer[10][0][3] [6]), .QN());
   DFF_X1 \buffer_reg[10][0][3][5]  (.D(\input_filter[0][3] [5]), .CK(n_56_7), 
      .Q(\buffer[10][0][3] [5]), .QN());
   DFF_X1 \buffer_reg[10][0][3][4]  (.D(\input_filter[0][3] [4]), .CK(n_56_7), 
      .Q(\buffer[10][0][3] [4]), .QN());
   DFF_X1 \buffer_reg[10][0][3][3]  (.D(\input_filter[0][3] [3]), .CK(n_56_7), 
      .Q(\buffer[10][0][3] [3]), .QN());
   DFF_X1 \buffer_reg[10][0][3][2]  (.D(\input_filter[0][3] [2]), .CK(n_56_7), 
      .Q(\buffer[10][0][3] [2]), .QN());
   DFF_X1 \buffer_reg[10][0][3][1]  (.D(\input_filter[0][3] [1]), .CK(n_56_7), 
      .Q(\buffer[10][0][3] [1]), .QN());
   DFF_X1 \buffer_reg[10][0][3][0]  (.D(\input_filter[0][3] [0]), .CK(n_56_7), 
      .Q(\buffer[10][0][3] [0]), .QN());
   DFF_X1 \buffer_reg[11][0][3][15]  (.D(\input_filter[0][3] [15]), .CK(n_56_8), 
      .Q(\buffer[11][0][3] [15]), .QN());
   DFF_X1 \buffer_reg[11][0][3][14]  (.D(\input_filter[0][3] [14]), .CK(n_56_8), 
      .Q(\buffer[11][0][3] [14]), .QN());
   DFF_X1 \buffer_reg[11][0][3][13]  (.D(\input_filter[0][3] [13]), .CK(n_56_8), 
      .Q(\buffer[11][0][3] [13]), .QN());
   DFF_X1 \buffer_reg[11][0][3][12]  (.D(\input_filter[0][3] [12]), .CK(n_56_8), 
      .Q(\buffer[11][0][3] [12]), .QN());
   DFF_X1 \buffer_reg[11][0][3][11]  (.D(\input_filter[0][3] [11]), .CK(n_56_8), 
      .Q(\buffer[11][0][3] [11]), .QN());
   DFF_X1 \buffer_reg[11][0][3][10]  (.D(\input_filter[0][3] [10]), .CK(n_56_8), 
      .Q(\buffer[11][0][3] [10]), .QN());
   DFF_X1 \buffer_reg[11][0][3][9]  (.D(\input_filter[0][3] [9]), .CK(n_56_8), 
      .Q(\buffer[11][0][3] [9]), .QN());
   DFF_X1 \buffer_reg[11][0][3][8]  (.D(\input_filter[0][3] [8]), .CK(n_56_8), 
      .Q(\buffer[11][0][3] [8]), .QN());
   DFF_X1 \buffer_reg[11][0][3][7]  (.D(\input_filter[0][3] [7]), .CK(n_56_8), 
      .Q(\buffer[11][0][3] [7]), .QN());
   DFF_X1 \buffer_reg[11][0][3][6]  (.D(\input_filter[0][3] [6]), .CK(n_56_8), 
      .Q(\buffer[11][0][3] [6]), .QN());
   DFF_X1 \buffer_reg[11][0][3][5]  (.D(\input_filter[0][3] [5]), .CK(n_56_8), 
      .Q(\buffer[11][0][3] [5]), .QN());
   DFF_X1 \buffer_reg[11][0][3][4]  (.D(\input_filter[0][3] [4]), .CK(n_56_8), 
      .Q(\buffer[11][0][3] [4]), .QN());
   DFF_X1 \buffer_reg[11][0][3][3]  (.D(\input_filter[0][3] [3]), .CK(n_56_8), 
      .Q(\buffer[11][0][3] [3]), .QN());
   DFF_X1 \buffer_reg[11][0][3][2]  (.D(\input_filter[0][3] [2]), .CK(n_56_8), 
      .Q(\buffer[11][0][3] [2]), .QN());
   DFF_X1 \buffer_reg[11][0][3][1]  (.D(\input_filter[0][3] [1]), .CK(n_56_8), 
      .Q(\buffer[11][0][3] [1]), .QN());
   DFF_X1 \buffer_reg[11][0][3][0]  (.D(\input_filter[0][3] [0]), .CK(n_56_8), 
      .Q(\buffer[11][0][3] [0]), .QN());
   DFF_X1 \buffer_reg[12][0][3][15]  (.D(\input_filter[0][3] [15]), .CK(n_56_9), 
      .Q(\buffer[12][0][3] [15]), .QN());
   DFF_X1 \buffer_reg[12][0][3][14]  (.D(\input_filter[0][3] [14]), .CK(n_56_9), 
      .Q(\buffer[12][0][3] [14]), .QN());
   DFF_X1 \buffer_reg[12][0][3][13]  (.D(\input_filter[0][3] [13]), .CK(n_56_9), 
      .Q(\buffer[12][0][3] [13]), .QN());
   DFF_X1 \buffer_reg[12][0][3][12]  (.D(\input_filter[0][3] [12]), .CK(n_56_9), 
      .Q(\buffer[12][0][3] [12]), .QN());
   DFF_X1 \buffer_reg[12][0][3][11]  (.D(\input_filter[0][3] [11]), .CK(n_56_9), 
      .Q(\buffer[12][0][3] [11]), .QN());
   DFF_X1 \buffer_reg[12][0][3][10]  (.D(\input_filter[0][3] [10]), .CK(n_56_9), 
      .Q(\buffer[12][0][3] [10]), .QN());
   DFF_X1 \buffer_reg[12][0][3][9]  (.D(\input_filter[0][3] [9]), .CK(n_56_9), 
      .Q(\buffer[12][0][3] [9]), .QN());
   DFF_X1 \buffer_reg[12][0][3][8]  (.D(\input_filter[0][3] [8]), .CK(n_56_9), 
      .Q(\buffer[12][0][3] [8]), .QN());
   DFF_X1 \buffer_reg[12][0][3][7]  (.D(\input_filter[0][3] [7]), .CK(n_56_9), 
      .Q(\buffer[12][0][3] [7]), .QN());
   DFF_X1 \buffer_reg[12][0][3][6]  (.D(\input_filter[0][3] [6]), .CK(n_56_9), 
      .Q(\buffer[12][0][3] [6]), .QN());
   DFF_X1 \buffer_reg[12][0][3][5]  (.D(\input_filter[0][3] [5]), .CK(n_56_9), 
      .Q(\buffer[12][0][3] [5]), .QN());
   DFF_X1 \buffer_reg[12][0][3][4]  (.D(\input_filter[0][3] [4]), .CK(n_56_9), 
      .Q(\buffer[12][0][3] [4]), .QN());
   DFF_X1 \buffer_reg[12][0][3][3]  (.D(\input_filter[0][3] [3]), .CK(n_56_9), 
      .Q(\buffer[12][0][3] [3]), .QN());
   DFF_X1 \buffer_reg[12][0][3][2]  (.D(\input_filter[0][3] [2]), .CK(n_56_9), 
      .Q(\buffer[12][0][3] [2]), .QN());
   DFF_X1 \buffer_reg[12][0][3][1]  (.D(\input_filter[0][3] [1]), .CK(n_56_9), 
      .Q(\buffer[12][0][3] [1]), .QN());
   DFF_X1 \buffer_reg[12][0][3][0]  (.D(\input_filter[0][3] [0]), .CK(n_56_9), 
      .Q(\buffer[12][0][3] [0]), .QN());
   DFF_X1 \buffer_reg[13][0][3][15]  (.D(\input_filter[0][3] [15]), .CK(n_56_10), 
      .Q(\buffer[13][0][3] [15]), .QN());
   DFF_X1 \buffer_reg[13][0][3][14]  (.D(\input_filter[0][3] [14]), .CK(n_56_10), 
      .Q(\buffer[13][0][3] [14]), .QN());
   DFF_X1 \buffer_reg[13][0][3][13]  (.D(\input_filter[0][3] [13]), .CK(n_56_10), 
      .Q(\buffer[13][0][3] [13]), .QN());
   DFF_X1 \buffer_reg[13][0][3][12]  (.D(\input_filter[0][3] [12]), .CK(n_56_10), 
      .Q(\buffer[13][0][3] [12]), .QN());
   DFF_X1 \buffer_reg[13][0][3][11]  (.D(\input_filter[0][3] [11]), .CK(n_56_10), 
      .Q(\buffer[13][0][3] [11]), .QN());
   DFF_X1 \buffer_reg[13][0][3][10]  (.D(\input_filter[0][3] [10]), .CK(n_56_10), 
      .Q(\buffer[13][0][3] [10]), .QN());
   DFF_X1 \buffer_reg[13][0][3][9]  (.D(\input_filter[0][3] [9]), .CK(n_56_10), 
      .Q(\buffer[13][0][3] [9]), .QN());
   DFF_X1 \buffer_reg[13][0][3][8]  (.D(\input_filter[0][3] [8]), .CK(n_56_10), 
      .Q(\buffer[13][0][3] [8]), .QN());
   DFF_X1 \buffer_reg[13][0][3][7]  (.D(\input_filter[0][3] [7]), .CK(n_56_10), 
      .Q(\buffer[13][0][3] [7]), .QN());
   DFF_X1 \buffer_reg[13][0][3][6]  (.D(\input_filter[0][3] [6]), .CK(n_56_10), 
      .Q(\buffer[13][0][3] [6]), .QN());
   DFF_X1 \buffer_reg[13][0][3][5]  (.D(\input_filter[0][3] [5]), .CK(n_56_10), 
      .Q(\buffer[13][0][3] [5]), .QN());
   DFF_X1 \buffer_reg[13][0][3][4]  (.D(\input_filter[0][3] [4]), .CK(n_56_10), 
      .Q(\buffer[13][0][3] [4]), .QN());
   DFF_X1 \buffer_reg[13][0][3][3]  (.D(\input_filter[0][3] [3]), .CK(n_56_10), 
      .Q(\buffer[13][0][3] [3]), .QN());
   DFF_X1 \buffer_reg[13][0][3][2]  (.D(\input_filter[0][3] [2]), .CK(n_56_10), 
      .Q(\buffer[13][0][3] [2]), .QN());
   DFF_X1 \buffer_reg[13][0][3][1]  (.D(\input_filter[0][3] [1]), .CK(n_56_10), 
      .Q(\buffer[13][0][3] [1]), .QN());
   DFF_X1 \buffer_reg[13][0][3][0]  (.D(\input_filter[0][3] [0]), .CK(n_56_10), 
      .Q(\buffer[13][0][3] [0]), .QN());
   DFF_X1 \buffer_reg[14][0][3][15]  (.D(\input_filter[0][3] [15]), .CK(n_56_11), 
      .Q(\buffer[14][0][3] [15]), .QN());
   DFF_X1 \buffer_reg[14][0][3][14]  (.D(\input_filter[0][3] [14]), .CK(n_56_11), 
      .Q(\buffer[14][0][3] [14]), .QN());
   DFF_X1 \buffer_reg[14][0][3][13]  (.D(\input_filter[0][3] [13]), .CK(n_56_11), 
      .Q(\buffer[14][0][3] [13]), .QN());
   DFF_X1 \buffer_reg[14][0][3][12]  (.D(\input_filter[0][3] [12]), .CK(n_56_11), 
      .Q(\buffer[14][0][3] [12]), .QN());
   DFF_X1 \buffer_reg[14][0][3][11]  (.D(\input_filter[0][3] [11]), .CK(n_56_11), 
      .Q(\buffer[14][0][3] [11]), .QN());
   DFF_X1 \buffer_reg[14][0][3][10]  (.D(\input_filter[0][3] [10]), .CK(n_56_11), 
      .Q(\buffer[14][0][3] [10]), .QN());
   DFF_X1 \buffer_reg[14][0][3][9]  (.D(\input_filter[0][3] [9]), .CK(n_56_11), 
      .Q(\buffer[14][0][3] [9]), .QN());
   DFF_X1 \buffer_reg[14][0][3][8]  (.D(\input_filter[0][3] [8]), .CK(n_56_11), 
      .Q(\buffer[14][0][3] [8]), .QN());
   DFF_X1 \buffer_reg[14][0][3][7]  (.D(\input_filter[0][3] [7]), .CK(n_56_11), 
      .Q(\buffer[14][0][3] [7]), .QN());
   DFF_X1 \buffer_reg[14][0][3][6]  (.D(\input_filter[0][3] [6]), .CK(n_56_11), 
      .Q(\buffer[14][0][3] [6]), .QN());
   DFF_X1 \buffer_reg[14][0][3][5]  (.D(\input_filter[0][3] [5]), .CK(n_56_11), 
      .Q(\buffer[14][0][3] [5]), .QN());
   DFF_X1 \buffer_reg[14][0][3][4]  (.D(\input_filter[0][3] [4]), .CK(n_56_11), 
      .Q(\buffer[14][0][3] [4]), .QN());
   DFF_X1 \buffer_reg[14][0][3][3]  (.D(\input_filter[0][3] [3]), .CK(n_56_11), 
      .Q(\buffer[14][0][3] [3]), .QN());
   DFF_X1 \buffer_reg[14][0][3][2]  (.D(\input_filter[0][3] [2]), .CK(n_56_11), 
      .Q(\buffer[14][0][3] [2]), .QN());
   DFF_X1 \buffer_reg[14][0][3][1]  (.D(\input_filter[0][3] [1]), .CK(n_56_11), 
      .Q(\buffer[14][0][3] [1]), .QN());
   DFF_X1 \buffer_reg[14][0][3][0]  (.D(\input_filter[0][3] [0]), .CK(n_56_11), 
      .Q(\buffer[14][0][3] [0]), .QN());
   DFF_X1 \buffer_reg[15][0][3][15]  (.D(\input_filter[0][3] [15]), .CK(n_56_15), 
      .Q(\buffer[15][0][3] [15]), .QN());
   DFF_X1 \buffer_reg[15][0][3][14]  (.D(\input_filter[0][3] [14]), .CK(n_56_15), 
      .Q(\buffer[15][0][3] [14]), .QN());
   DFF_X1 \buffer_reg[15][0][3][13]  (.D(\input_filter[0][3] [13]), .CK(n_56_15), 
      .Q(\buffer[15][0][3] [13]), .QN());
   DFF_X1 \buffer_reg[15][0][3][12]  (.D(\input_filter[0][3] [12]), .CK(n_56_15), 
      .Q(\buffer[15][0][3] [12]), .QN());
   DFF_X1 \buffer_reg[15][0][3][11]  (.D(\input_filter[0][3] [11]), .CK(n_56_15), 
      .Q(\buffer[15][0][3] [11]), .QN());
   DFF_X1 \buffer_reg[15][0][3][10]  (.D(\input_filter[0][3] [10]), .CK(n_56_15), 
      .Q(\buffer[15][0][3] [10]), .QN());
   DFF_X1 \buffer_reg[15][0][3][9]  (.D(\input_filter[0][3] [9]), .CK(n_56_15), 
      .Q(\buffer[15][0][3] [9]), .QN());
   DFF_X1 \buffer_reg[15][0][3][8]  (.D(\input_filter[0][3] [8]), .CK(n_56_15), 
      .Q(\buffer[15][0][3] [8]), .QN());
   DFF_X1 \buffer_reg[15][0][3][7]  (.D(\input_filter[0][3] [7]), .CK(n_56_15), 
      .Q(\buffer[15][0][3] [7]), .QN());
   DFF_X1 \buffer_reg[15][0][3][6]  (.D(\input_filter[0][3] [6]), .CK(n_56_15), 
      .Q(\buffer[15][0][3] [6]), .QN());
   DFF_X1 \buffer_reg[15][0][3][5]  (.D(\input_filter[0][3] [5]), .CK(n_56_15), 
      .Q(\buffer[15][0][3] [5]), .QN());
   DFF_X1 \buffer_reg[15][0][3][4]  (.D(\input_filter[0][3] [4]), .CK(n_56_15), 
      .Q(\buffer[15][0][3] [4]), .QN());
   DFF_X1 \buffer_reg[15][0][3][3]  (.D(\input_filter[0][3] [3]), .CK(n_56_15), 
      .Q(\buffer[15][0][3] [3]), .QN());
   DFF_X1 \buffer_reg[15][0][3][2]  (.D(\input_filter[0][3] [2]), .CK(n_56_15), 
      .Q(\buffer[15][0][3] [2]), .QN());
   DFF_X1 \buffer_reg[15][0][3][1]  (.D(\input_filter[0][3] [1]), .CK(n_56_15), 
      .Q(\buffer[15][0][3] [1]), .QN());
   DFF_X1 \buffer_reg[15][0][3][0]  (.D(\input_filter[0][3] [0]), .CK(n_56_15), 
      .Q(\buffer[15][0][3] [0]), .QN());
   DFF_X1 \buffer_reg[0][1][0][15]  (.D(\input_filter[1][0] [15]), .CK(n_56_12), 
      .Q(\buffer[0][1][0] [15]), .QN());
   DFF_X1 \buffer_reg[0][1][0][14]  (.D(\input_filter[1][0] [14]), .CK(n_56_12), 
      .Q(\buffer[0][1][0] [14]), .QN());
   DFF_X1 \buffer_reg[0][1][0][13]  (.D(\input_filter[1][0] [13]), .CK(n_56_12), 
      .Q(\buffer[0][1][0] [13]), .QN());
   DFF_X1 \buffer_reg[0][1][0][12]  (.D(\input_filter[1][0] [12]), .CK(n_56_12), 
      .Q(\buffer[0][1][0] [12]), .QN());
   DFF_X1 \buffer_reg[0][1][0][11]  (.D(\input_filter[1][0] [11]), .CK(n_56_12), 
      .Q(\buffer[0][1][0] [11]), .QN());
   DFF_X1 \buffer_reg[0][1][0][10]  (.D(\input_filter[1][0] [10]), .CK(n_56_12), 
      .Q(\buffer[0][1][0] [10]), .QN());
   DFF_X1 \buffer_reg[0][1][0][9]  (.D(\input_filter[1][0] [9]), .CK(n_56_12), 
      .Q(\buffer[0][1][0] [9]), .QN());
   DFF_X1 \buffer_reg[0][1][0][8]  (.D(\input_filter[1][0] [8]), .CK(n_56_12), 
      .Q(\buffer[0][1][0] [8]), .QN());
   DFF_X1 \buffer_reg[0][1][0][7]  (.D(\input_filter[1][0] [7]), .CK(n_56_12), 
      .Q(\buffer[0][1][0] [7]), .QN());
   DFF_X1 \buffer_reg[0][1][0][6]  (.D(\input_filter[1][0] [6]), .CK(n_56_12), 
      .Q(\buffer[0][1][0] [6]), .QN());
   DFF_X1 \buffer_reg[0][1][0][5]  (.D(\input_filter[1][0] [5]), .CK(n_56_12), 
      .Q(\buffer[0][1][0] [5]), .QN());
   DFF_X1 \buffer_reg[0][1][0][4]  (.D(\input_filter[1][0] [4]), .CK(n_56_12), 
      .Q(\buffer[0][1][0] [4]), .QN());
   DFF_X1 \buffer_reg[0][1][0][3]  (.D(\input_filter[1][0] [3]), .CK(n_56_12), 
      .Q(\buffer[0][1][0] [3]), .QN());
   DFF_X1 \buffer_reg[0][1][0][2]  (.D(\input_filter[1][0] [2]), .CK(n_56_12), 
      .Q(\buffer[0][1][0] [2]), .QN());
   DFF_X1 \buffer_reg[0][1][0][1]  (.D(\input_filter[1][0] [1]), .CK(n_56_12), 
      .Q(\buffer[0][1][0] [1]), .QN());
   DFF_X1 \buffer_reg[0][1][0][0]  (.D(\input_filter[1][0] [0]), .CK(n_56_12), 
      .Q(\buffer[0][1][0] [0]), .QN());
   DFF_X1 \buffer_reg[1][1][0][15]  (.D(\input_filter[1][0] [15]), .CK(n_56_13), 
      .Q(\buffer[1][1][0] [15]), .QN());
   DFF_X1 \buffer_reg[1][1][0][14]  (.D(\input_filter[1][0] [14]), .CK(n_56_13), 
      .Q(\buffer[1][1][0] [14]), .QN());
   DFF_X1 \buffer_reg[1][1][0][13]  (.D(\input_filter[1][0] [13]), .CK(n_56_13), 
      .Q(\buffer[1][1][0] [13]), .QN());
   DFF_X1 \buffer_reg[1][1][0][12]  (.D(\input_filter[1][0] [12]), .CK(n_56_13), 
      .Q(\buffer[1][1][0] [12]), .QN());
   DFF_X1 \buffer_reg[1][1][0][11]  (.D(\input_filter[1][0] [11]), .CK(n_56_13), 
      .Q(\buffer[1][1][0] [11]), .QN());
   DFF_X1 \buffer_reg[1][1][0][10]  (.D(\input_filter[1][0] [10]), .CK(n_56_13), 
      .Q(\buffer[1][1][0] [10]), .QN());
   DFF_X1 \buffer_reg[1][1][0][9]  (.D(\input_filter[1][0] [9]), .CK(n_56_13), 
      .Q(\buffer[1][1][0] [9]), .QN());
   DFF_X1 \buffer_reg[1][1][0][8]  (.D(\input_filter[1][0] [8]), .CK(n_56_13), 
      .Q(\buffer[1][1][0] [8]), .QN());
   DFF_X1 \buffer_reg[1][1][0][7]  (.D(\input_filter[1][0] [7]), .CK(n_56_13), 
      .Q(\buffer[1][1][0] [7]), .QN());
   DFF_X1 \buffer_reg[1][1][0][6]  (.D(\input_filter[1][0] [6]), .CK(n_56_13), 
      .Q(\buffer[1][1][0] [6]), .QN());
   DFF_X1 \buffer_reg[1][1][0][5]  (.D(\input_filter[1][0] [5]), .CK(n_56_13), 
      .Q(\buffer[1][1][0] [5]), .QN());
   DFF_X1 \buffer_reg[1][1][0][4]  (.D(\input_filter[1][0] [4]), .CK(n_56_13), 
      .Q(\buffer[1][1][0] [4]), .QN());
   DFF_X1 \buffer_reg[1][1][0][3]  (.D(\input_filter[1][0] [3]), .CK(n_56_13), 
      .Q(\buffer[1][1][0] [3]), .QN());
   DFF_X1 \buffer_reg[1][1][0][2]  (.D(\input_filter[1][0] [2]), .CK(n_56_13), 
      .Q(\buffer[1][1][0] [2]), .QN());
   DFF_X1 \buffer_reg[1][1][0][1]  (.D(\input_filter[1][0] [1]), .CK(n_56_13), 
      .Q(\buffer[1][1][0] [1]), .QN());
   DFF_X1 \buffer_reg[1][1][0][0]  (.D(\input_filter[1][0] [0]), .CK(n_56_13), 
      .Q(\buffer[1][1][0] [0]), .QN());
   DFF_X1 \buffer_reg[2][1][0][15]  (.D(\input_filter[1][0] [15]), .CK(n_56_14), 
      .Q(\buffer[2][1][0] [15]), .QN());
   DFF_X1 \buffer_reg[2][1][0][14]  (.D(\input_filter[1][0] [14]), .CK(n_56_14), 
      .Q(\buffer[2][1][0] [14]), .QN());
   DFF_X1 \buffer_reg[2][1][0][13]  (.D(\input_filter[1][0] [13]), .CK(n_56_14), 
      .Q(\buffer[2][1][0] [13]), .QN());
   DFF_X1 \buffer_reg[2][1][0][12]  (.D(\input_filter[1][0] [12]), .CK(n_56_14), 
      .Q(\buffer[2][1][0] [12]), .QN());
   DFF_X1 \buffer_reg[2][1][0][11]  (.D(\input_filter[1][0] [11]), .CK(n_56_14), 
      .Q(\buffer[2][1][0] [11]), .QN());
   DFF_X1 \buffer_reg[2][1][0][10]  (.D(\input_filter[1][0] [10]), .CK(n_56_14), 
      .Q(\buffer[2][1][0] [10]), .QN());
   DFF_X1 \buffer_reg[2][1][0][9]  (.D(\input_filter[1][0] [9]), .CK(n_56_14), 
      .Q(\buffer[2][1][0] [9]), .QN());
   DFF_X1 \buffer_reg[2][1][0][8]  (.D(\input_filter[1][0] [8]), .CK(n_56_14), 
      .Q(\buffer[2][1][0] [8]), .QN());
   DFF_X1 \buffer_reg[2][1][0][7]  (.D(\input_filter[1][0] [7]), .CK(n_56_14), 
      .Q(\buffer[2][1][0] [7]), .QN());
   DFF_X1 \buffer_reg[2][1][0][6]  (.D(\input_filter[1][0] [6]), .CK(n_56_14), 
      .Q(\buffer[2][1][0] [6]), .QN());
   DFF_X1 \buffer_reg[2][1][0][5]  (.D(\input_filter[1][0] [5]), .CK(n_56_14), 
      .Q(\buffer[2][1][0] [5]), .QN());
   DFF_X1 \buffer_reg[2][1][0][4]  (.D(\input_filter[1][0] [4]), .CK(n_56_14), 
      .Q(\buffer[2][1][0] [4]), .QN());
   DFF_X1 \buffer_reg[2][1][0][3]  (.D(\input_filter[1][0] [3]), .CK(n_56_14), 
      .Q(\buffer[2][1][0] [3]), .QN());
   DFF_X1 \buffer_reg[2][1][0][2]  (.D(\input_filter[1][0] [2]), .CK(n_56_14), 
      .Q(\buffer[2][1][0] [2]), .QN());
   DFF_X1 \buffer_reg[2][1][0][1]  (.D(\input_filter[1][0] [1]), .CK(n_56_14), 
      .Q(\buffer[2][1][0] [1]), .QN());
   DFF_X1 \buffer_reg[2][1][0][0]  (.D(\input_filter[1][0] [0]), .CK(n_56_14), 
      .Q(\buffer[2][1][0] [0]), .QN());
   DFF_X1 \buffer_reg[3][1][0][15]  (.D(\input_filter[1][0] [15]), .CK(n_56_0), 
      .Q(\buffer[3][1][0] [15]), .QN());
   DFF_X1 \buffer_reg[3][1][0][14]  (.D(\input_filter[1][0] [14]), .CK(n_56_0), 
      .Q(\buffer[3][1][0] [14]), .QN());
   DFF_X1 \buffer_reg[3][1][0][13]  (.D(\input_filter[1][0] [13]), .CK(n_56_0), 
      .Q(\buffer[3][1][0] [13]), .QN());
   DFF_X1 \buffer_reg[3][1][0][12]  (.D(\input_filter[1][0] [12]), .CK(n_56_0), 
      .Q(\buffer[3][1][0] [12]), .QN());
   DFF_X1 \buffer_reg[3][1][0][11]  (.D(\input_filter[1][0] [11]), .CK(n_56_0), 
      .Q(\buffer[3][1][0] [11]), .QN());
   DFF_X1 \buffer_reg[3][1][0][10]  (.D(\input_filter[1][0] [10]), .CK(n_56_0), 
      .Q(\buffer[3][1][0] [10]), .QN());
   DFF_X1 \buffer_reg[3][1][0][9]  (.D(\input_filter[1][0] [9]), .CK(n_56_0), 
      .Q(\buffer[3][1][0] [9]), .QN());
   DFF_X1 \buffer_reg[3][1][0][8]  (.D(\input_filter[1][0] [8]), .CK(n_56_0), 
      .Q(\buffer[3][1][0] [8]), .QN());
   DFF_X1 \buffer_reg[3][1][0][7]  (.D(\input_filter[1][0] [7]), .CK(n_56_0), 
      .Q(\buffer[3][1][0] [7]), .QN());
   DFF_X1 \buffer_reg[3][1][0][6]  (.D(\input_filter[1][0] [6]), .CK(n_56_0), 
      .Q(\buffer[3][1][0] [6]), .QN());
   DFF_X1 \buffer_reg[3][1][0][5]  (.D(\input_filter[1][0] [5]), .CK(n_56_0), 
      .Q(\buffer[3][1][0] [5]), .QN());
   DFF_X1 \buffer_reg[3][1][0][4]  (.D(\input_filter[1][0] [4]), .CK(n_56_0), 
      .Q(\buffer[3][1][0] [4]), .QN());
   DFF_X1 \buffer_reg[3][1][0][3]  (.D(\input_filter[1][0] [3]), .CK(n_56_0), 
      .Q(\buffer[3][1][0] [3]), .QN());
   DFF_X1 \buffer_reg[3][1][0][2]  (.D(\input_filter[1][0] [2]), .CK(n_56_0), 
      .Q(\buffer[3][1][0] [2]), .QN());
   DFF_X1 \buffer_reg[3][1][0][1]  (.D(\input_filter[1][0] [1]), .CK(n_56_0), 
      .Q(\buffer[3][1][0] [1]), .QN());
   DFF_X1 \buffer_reg[3][1][0][0]  (.D(\input_filter[1][0] [0]), .CK(n_56_0), 
      .Q(\buffer[3][1][0] [0]), .QN());
   DFF_X1 \buffer_reg[4][1][0][15]  (.D(\input_filter[1][0] [15]), .CK(n_56_1), 
      .Q(\buffer[4][1][0] [15]), .QN());
   DFF_X1 \buffer_reg[4][1][0][14]  (.D(\input_filter[1][0] [14]), .CK(n_56_1), 
      .Q(\buffer[4][1][0] [14]), .QN());
   DFF_X1 \buffer_reg[4][1][0][13]  (.D(\input_filter[1][0] [13]), .CK(n_56_1), 
      .Q(\buffer[4][1][0] [13]), .QN());
   DFF_X1 \buffer_reg[4][1][0][12]  (.D(\input_filter[1][0] [12]), .CK(n_56_1), 
      .Q(\buffer[4][1][0] [12]), .QN());
   DFF_X1 \buffer_reg[4][1][0][11]  (.D(\input_filter[1][0] [11]), .CK(n_56_1), 
      .Q(\buffer[4][1][0] [11]), .QN());
   DFF_X1 \buffer_reg[4][1][0][10]  (.D(\input_filter[1][0] [10]), .CK(n_56_1), 
      .Q(\buffer[4][1][0] [10]), .QN());
   DFF_X1 \buffer_reg[4][1][0][9]  (.D(\input_filter[1][0] [9]), .CK(n_56_1), 
      .Q(\buffer[4][1][0] [9]), .QN());
   DFF_X1 \buffer_reg[4][1][0][8]  (.D(\input_filter[1][0] [8]), .CK(n_56_1), 
      .Q(\buffer[4][1][0] [8]), .QN());
   DFF_X1 \buffer_reg[4][1][0][7]  (.D(\input_filter[1][0] [7]), .CK(n_56_1), 
      .Q(\buffer[4][1][0] [7]), .QN());
   DFF_X1 \buffer_reg[4][1][0][6]  (.D(\input_filter[1][0] [6]), .CK(n_56_1), 
      .Q(\buffer[4][1][0] [6]), .QN());
   DFF_X1 \buffer_reg[4][1][0][5]  (.D(\input_filter[1][0] [5]), .CK(n_56_1), 
      .Q(\buffer[4][1][0] [5]), .QN());
   DFF_X1 \buffer_reg[4][1][0][4]  (.D(\input_filter[1][0] [4]), .CK(n_56_1), 
      .Q(\buffer[4][1][0] [4]), .QN());
   DFF_X1 \buffer_reg[4][1][0][3]  (.D(\input_filter[1][0] [3]), .CK(n_56_1), 
      .Q(\buffer[4][1][0] [3]), .QN());
   DFF_X1 \buffer_reg[4][1][0][2]  (.D(\input_filter[1][0] [2]), .CK(n_56_1), 
      .Q(\buffer[4][1][0] [2]), .QN());
   DFF_X1 \buffer_reg[4][1][0][1]  (.D(\input_filter[1][0] [1]), .CK(n_56_1), 
      .Q(\buffer[4][1][0] [1]), .QN());
   DFF_X1 \buffer_reg[4][1][0][0]  (.D(\input_filter[1][0] [0]), .CK(n_56_1), 
      .Q(\buffer[4][1][0] [0]), .QN());
   DFF_X1 \buffer_reg[5][1][0][15]  (.D(\input_filter[1][0] [15]), .CK(n_56_2), 
      .Q(\buffer[5][1][0] [15]), .QN());
   DFF_X1 \buffer_reg[5][1][0][14]  (.D(\input_filter[1][0] [14]), .CK(n_56_2), 
      .Q(\buffer[5][1][0] [14]), .QN());
   DFF_X1 \buffer_reg[5][1][0][13]  (.D(\input_filter[1][0] [13]), .CK(n_56_2), 
      .Q(\buffer[5][1][0] [13]), .QN());
   DFF_X1 \buffer_reg[5][1][0][12]  (.D(\input_filter[1][0] [12]), .CK(n_56_2), 
      .Q(\buffer[5][1][0] [12]), .QN());
   DFF_X1 \buffer_reg[5][1][0][11]  (.D(\input_filter[1][0] [11]), .CK(n_56_2), 
      .Q(\buffer[5][1][0] [11]), .QN());
   DFF_X1 \buffer_reg[5][1][0][10]  (.D(\input_filter[1][0] [10]), .CK(n_56_2), 
      .Q(\buffer[5][1][0] [10]), .QN());
   DFF_X1 \buffer_reg[5][1][0][9]  (.D(\input_filter[1][0] [9]), .CK(n_56_2), 
      .Q(\buffer[5][1][0] [9]), .QN());
   DFF_X1 \buffer_reg[5][1][0][8]  (.D(\input_filter[1][0] [8]), .CK(n_56_2), 
      .Q(\buffer[5][1][0] [8]), .QN());
   DFF_X1 \buffer_reg[5][1][0][7]  (.D(\input_filter[1][0] [7]), .CK(n_56_2), 
      .Q(\buffer[5][1][0] [7]), .QN());
   DFF_X1 \buffer_reg[5][1][0][6]  (.D(\input_filter[1][0] [6]), .CK(n_56_2), 
      .Q(\buffer[5][1][0] [6]), .QN());
   DFF_X1 \buffer_reg[5][1][0][5]  (.D(\input_filter[1][0] [5]), .CK(n_56_2), 
      .Q(\buffer[5][1][0] [5]), .QN());
   DFF_X1 \buffer_reg[5][1][0][4]  (.D(\input_filter[1][0] [4]), .CK(n_56_2), 
      .Q(\buffer[5][1][0] [4]), .QN());
   DFF_X1 \buffer_reg[5][1][0][3]  (.D(\input_filter[1][0] [3]), .CK(n_56_2), 
      .Q(\buffer[5][1][0] [3]), .QN());
   DFF_X1 \buffer_reg[5][1][0][2]  (.D(\input_filter[1][0] [2]), .CK(n_56_2), 
      .Q(\buffer[5][1][0] [2]), .QN());
   DFF_X1 \buffer_reg[5][1][0][1]  (.D(\input_filter[1][0] [1]), .CK(n_56_2), 
      .Q(\buffer[5][1][0] [1]), .QN());
   DFF_X1 \buffer_reg[5][1][0][0]  (.D(\input_filter[1][0] [0]), .CK(n_56_2), 
      .Q(\buffer[5][1][0] [0]), .QN());
   DFF_X1 \buffer_reg[6][1][0][15]  (.D(\input_filter[1][0] [15]), .CK(n_56_3), 
      .Q(\buffer[6][1][0] [15]), .QN());
   DFF_X1 \buffer_reg[6][1][0][14]  (.D(\input_filter[1][0] [14]), .CK(n_56_3), 
      .Q(\buffer[6][1][0] [14]), .QN());
   DFF_X1 \buffer_reg[6][1][0][13]  (.D(\input_filter[1][0] [13]), .CK(n_56_3), 
      .Q(\buffer[6][1][0] [13]), .QN());
   DFF_X1 \buffer_reg[6][1][0][12]  (.D(\input_filter[1][0] [12]), .CK(n_56_3), 
      .Q(\buffer[6][1][0] [12]), .QN());
   DFF_X1 \buffer_reg[6][1][0][11]  (.D(\input_filter[1][0] [11]), .CK(n_56_3), 
      .Q(\buffer[6][1][0] [11]), .QN());
   DFF_X1 \buffer_reg[6][1][0][10]  (.D(\input_filter[1][0] [10]), .CK(n_56_3), 
      .Q(\buffer[6][1][0] [10]), .QN());
   DFF_X1 \buffer_reg[6][1][0][9]  (.D(\input_filter[1][0] [9]), .CK(n_56_3), 
      .Q(\buffer[6][1][0] [9]), .QN());
   DFF_X1 \buffer_reg[6][1][0][8]  (.D(\input_filter[1][0] [8]), .CK(n_56_3), 
      .Q(\buffer[6][1][0] [8]), .QN());
   DFF_X1 \buffer_reg[6][1][0][7]  (.D(\input_filter[1][0] [7]), .CK(n_56_3), 
      .Q(\buffer[6][1][0] [7]), .QN());
   DFF_X1 \buffer_reg[6][1][0][6]  (.D(\input_filter[1][0] [6]), .CK(n_56_3), 
      .Q(\buffer[6][1][0] [6]), .QN());
   DFF_X1 \buffer_reg[6][1][0][5]  (.D(\input_filter[1][0] [5]), .CK(n_56_3), 
      .Q(\buffer[6][1][0] [5]), .QN());
   DFF_X1 \buffer_reg[6][1][0][4]  (.D(\input_filter[1][0] [4]), .CK(n_56_3), 
      .Q(\buffer[6][1][0] [4]), .QN());
   DFF_X1 \buffer_reg[6][1][0][3]  (.D(\input_filter[1][0] [3]), .CK(n_56_3), 
      .Q(\buffer[6][1][0] [3]), .QN());
   DFF_X1 \buffer_reg[6][1][0][2]  (.D(\input_filter[1][0] [2]), .CK(n_56_3), 
      .Q(\buffer[6][1][0] [2]), .QN());
   DFF_X1 \buffer_reg[6][1][0][1]  (.D(\input_filter[1][0] [1]), .CK(n_56_3), 
      .Q(\buffer[6][1][0] [1]), .QN());
   DFF_X1 \buffer_reg[6][1][0][0]  (.D(\input_filter[1][0] [0]), .CK(n_56_3), 
      .Q(\buffer[6][1][0] [0]), .QN());
   DFF_X1 \buffer_reg[7][1][0][15]  (.D(\input_filter[1][0] [15]), .CK(n_56_4), 
      .Q(\buffer[7][1][0] [15]), .QN());
   DFF_X1 \buffer_reg[7][1][0][14]  (.D(\input_filter[1][0] [14]), .CK(n_56_4), 
      .Q(\buffer[7][1][0] [14]), .QN());
   DFF_X1 \buffer_reg[7][1][0][13]  (.D(\input_filter[1][0] [13]), .CK(n_56_4), 
      .Q(\buffer[7][1][0] [13]), .QN());
   DFF_X1 \buffer_reg[7][1][0][12]  (.D(\input_filter[1][0] [12]), .CK(n_56_4), 
      .Q(\buffer[7][1][0] [12]), .QN());
   DFF_X1 \buffer_reg[7][1][0][11]  (.D(\input_filter[1][0] [11]), .CK(n_56_4), 
      .Q(\buffer[7][1][0] [11]), .QN());
   DFF_X1 \buffer_reg[7][1][0][10]  (.D(\input_filter[1][0] [10]), .CK(n_56_4), 
      .Q(\buffer[7][1][0] [10]), .QN());
   DFF_X1 \buffer_reg[7][1][0][9]  (.D(\input_filter[1][0] [9]), .CK(n_56_4), 
      .Q(\buffer[7][1][0] [9]), .QN());
   DFF_X1 \buffer_reg[7][1][0][8]  (.D(\input_filter[1][0] [8]), .CK(n_56_4), 
      .Q(\buffer[7][1][0] [8]), .QN());
   DFF_X1 \buffer_reg[7][1][0][7]  (.D(\input_filter[1][0] [7]), .CK(n_56_4), 
      .Q(\buffer[7][1][0] [7]), .QN());
   DFF_X1 \buffer_reg[7][1][0][6]  (.D(\input_filter[1][0] [6]), .CK(n_56_4), 
      .Q(\buffer[7][1][0] [6]), .QN());
   DFF_X1 \buffer_reg[7][1][0][5]  (.D(\input_filter[1][0] [5]), .CK(n_56_4), 
      .Q(\buffer[7][1][0] [5]), .QN());
   DFF_X1 \buffer_reg[7][1][0][4]  (.D(\input_filter[1][0] [4]), .CK(n_56_4), 
      .Q(\buffer[7][1][0] [4]), .QN());
   DFF_X1 \buffer_reg[7][1][0][3]  (.D(\input_filter[1][0] [3]), .CK(n_56_4), 
      .Q(\buffer[7][1][0] [3]), .QN());
   DFF_X1 \buffer_reg[7][1][0][2]  (.D(\input_filter[1][0] [2]), .CK(n_56_4), 
      .Q(\buffer[7][1][0] [2]), .QN());
   DFF_X1 \buffer_reg[7][1][0][1]  (.D(\input_filter[1][0] [1]), .CK(n_56_4), 
      .Q(\buffer[7][1][0] [1]), .QN());
   DFF_X1 \buffer_reg[7][1][0][0]  (.D(\input_filter[1][0] [0]), .CK(n_56_4), 
      .Q(\buffer[7][1][0] [0]), .QN());
   DFF_X1 \buffer_reg[8][1][0][15]  (.D(\input_filter[1][0] [15]), .CK(n_56_5), 
      .Q(\buffer[8][1][0] [15]), .QN());
   DFF_X1 \buffer_reg[8][1][0][14]  (.D(\input_filter[1][0] [14]), .CK(n_56_5), 
      .Q(\buffer[8][1][0] [14]), .QN());
   DFF_X1 \buffer_reg[8][1][0][13]  (.D(\input_filter[1][0] [13]), .CK(n_56_5), 
      .Q(\buffer[8][1][0] [13]), .QN());
   DFF_X1 \buffer_reg[8][1][0][12]  (.D(\input_filter[1][0] [12]), .CK(n_56_5), 
      .Q(\buffer[8][1][0] [12]), .QN());
   DFF_X1 \buffer_reg[8][1][0][11]  (.D(\input_filter[1][0] [11]), .CK(n_56_5), 
      .Q(\buffer[8][1][0] [11]), .QN());
   DFF_X1 \buffer_reg[8][1][0][10]  (.D(\input_filter[1][0] [10]), .CK(n_56_5), 
      .Q(\buffer[8][1][0] [10]), .QN());
   DFF_X1 \buffer_reg[8][1][0][9]  (.D(\input_filter[1][0] [9]), .CK(n_56_5), 
      .Q(\buffer[8][1][0] [9]), .QN());
   DFF_X1 \buffer_reg[8][1][0][8]  (.D(\input_filter[1][0] [8]), .CK(n_56_5), 
      .Q(\buffer[8][1][0] [8]), .QN());
   DFF_X1 \buffer_reg[8][1][0][7]  (.D(\input_filter[1][0] [7]), .CK(n_56_5), 
      .Q(\buffer[8][1][0] [7]), .QN());
   DFF_X1 \buffer_reg[8][1][0][6]  (.D(\input_filter[1][0] [6]), .CK(n_56_5), 
      .Q(\buffer[8][1][0] [6]), .QN());
   DFF_X1 \buffer_reg[8][1][0][5]  (.D(\input_filter[1][0] [5]), .CK(n_56_5), 
      .Q(\buffer[8][1][0] [5]), .QN());
   DFF_X1 \buffer_reg[8][1][0][4]  (.D(\input_filter[1][0] [4]), .CK(n_56_5), 
      .Q(\buffer[8][1][0] [4]), .QN());
   DFF_X1 \buffer_reg[8][1][0][3]  (.D(\input_filter[1][0] [3]), .CK(n_56_5), 
      .Q(\buffer[8][1][0] [3]), .QN());
   DFF_X1 \buffer_reg[8][1][0][2]  (.D(\input_filter[1][0] [2]), .CK(n_56_5), 
      .Q(\buffer[8][1][0] [2]), .QN());
   DFF_X1 \buffer_reg[8][1][0][1]  (.D(\input_filter[1][0] [1]), .CK(n_56_5), 
      .Q(\buffer[8][1][0] [1]), .QN());
   DFF_X1 \buffer_reg[8][1][0][0]  (.D(\input_filter[1][0] [0]), .CK(n_56_5), 
      .Q(\buffer[8][1][0] [0]), .QN());
   DFF_X1 \buffer_reg[9][1][0][15]  (.D(\input_filter[1][0] [15]), .CK(n_56_6), 
      .Q(\buffer[9][1][0] [15]), .QN());
   DFF_X1 \buffer_reg[9][1][0][14]  (.D(\input_filter[1][0] [14]), .CK(n_56_6), 
      .Q(\buffer[9][1][0] [14]), .QN());
   DFF_X1 \buffer_reg[9][1][0][13]  (.D(\input_filter[1][0] [13]), .CK(n_56_6), 
      .Q(\buffer[9][1][0] [13]), .QN());
   DFF_X1 \buffer_reg[9][1][0][12]  (.D(\input_filter[1][0] [12]), .CK(n_56_6), 
      .Q(\buffer[9][1][0] [12]), .QN());
   DFF_X1 \buffer_reg[9][1][0][11]  (.D(\input_filter[1][0] [11]), .CK(n_56_6), 
      .Q(\buffer[9][1][0] [11]), .QN());
   DFF_X1 \buffer_reg[9][1][0][10]  (.D(\input_filter[1][0] [10]), .CK(n_56_6), 
      .Q(\buffer[9][1][0] [10]), .QN());
   DFF_X1 \buffer_reg[9][1][0][9]  (.D(\input_filter[1][0] [9]), .CK(n_56_6), 
      .Q(\buffer[9][1][0] [9]), .QN());
   DFF_X1 \buffer_reg[9][1][0][8]  (.D(\input_filter[1][0] [8]), .CK(n_56_6), 
      .Q(\buffer[9][1][0] [8]), .QN());
   DFF_X1 \buffer_reg[9][1][0][7]  (.D(\input_filter[1][0] [7]), .CK(n_56_6), 
      .Q(\buffer[9][1][0] [7]), .QN());
   DFF_X1 \buffer_reg[9][1][0][6]  (.D(\input_filter[1][0] [6]), .CK(n_56_6), 
      .Q(\buffer[9][1][0] [6]), .QN());
   DFF_X1 \buffer_reg[9][1][0][5]  (.D(\input_filter[1][0] [5]), .CK(n_56_6), 
      .Q(\buffer[9][1][0] [5]), .QN());
   DFF_X1 \buffer_reg[9][1][0][4]  (.D(\input_filter[1][0] [4]), .CK(n_56_6), 
      .Q(\buffer[9][1][0] [4]), .QN());
   DFF_X1 \buffer_reg[9][1][0][3]  (.D(\input_filter[1][0] [3]), .CK(n_56_6), 
      .Q(\buffer[9][1][0] [3]), .QN());
   DFF_X1 \buffer_reg[9][1][0][2]  (.D(\input_filter[1][0] [2]), .CK(n_56_6), 
      .Q(\buffer[9][1][0] [2]), .QN());
   DFF_X1 \buffer_reg[9][1][0][1]  (.D(\input_filter[1][0] [1]), .CK(n_56_6), 
      .Q(\buffer[9][1][0] [1]), .QN());
   DFF_X1 \buffer_reg[9][1][0][0]  (.D(\input_filter[1][0] [0]), .CK(n_56_6), 
      .Q(\buffer[9][1][0] [0]), .QN());
   DFF_X1 \buffer_reg[10][1][0][15]  (.D(\input_filter[1][0] [15]), .CK(n_56_7), 
      .Q(\buffer[10][1][0] [15]), .QN());
   DFF_X1 \buffer_reg[10][1][0][14]  (.D(\input_filter[1][0] [14]), .CK(n_56_7), 
      .Q(\buffer[10][1][0] [14]), .QN());
   DFF_X1 \buffer_reg[10][1][0][13]  (.D(\input_filter[1][0] [13]), .CK(n_56_7), 
      .Q(\buffer[10][1][0] [13]), .QN());
   DFF_X1 \buffer_reg[10][1][0][12]  (.D(\input_filter[1][0] [12]), .CK(n_56_7), 
      .Q(\buffer[10][1][0] [12]), .QN());
   DFF_X1 \buffer_reg[10][1][0][11]  (.D(\input_filter[1][0] [11]), .CK(n_56_7), 
      .Q(\buffer[10][1][0] [11]), .QN());
   DFF_X1 \buffer_reg[10][1][0][10]  (.D(\input_filter[1][0] [10]), .CK(n_56_7), 
      .Q(\buffer[10][1][0] [10]), .QN());
   DFF_X1 \buffer_reg[10][1][0][9]  (.D(\input_filter[1][0] [9]), .CK(n_56_7), 
      .Q(\buffer[10][1][0] [9]), .QN());
   DFF_X1 \buffer_reg[10][1][0][8]  (.D(\input_filter[1][0] [8]), .CK(n_56_7), 
      .Q(\buffer[10][1][0] [8]), .QN());
   DFF_X1 \buffer_reg[10][1][0][7]  (.D(\input_filter[1][0] [7]), .CK(n_56_7), 
      .Q(\buffer[10][1][0] [7]), .QN());
   DFF_X1 \buffer_reg[10][1][0][6]  (.D(\input_filter[1][0] [6]), .CK(n_56_7), 
      .Q(\buffer[10][1][0] [6]), .QN());
   DFF_X1 \buffer_reg[10][1][0][5]  (.D(\input_filter[1][0] [5]), .CK(n_56_7), 
      .Q(\buffer[10][1][0] [5]), .QN());
   DFF_X1 \buffer_reg[10][1][0][4]  (.D(\input_filter[1][0] [4]), .CK(n_56_7), 
      .Q(\buffer[10][1][0] [4]), .QN());
   DFF_X1 \buffer_reg[10][1][0][3]  (.D(\input_filter[1][0] [3]), .CK(n_56_7), 
      .Q(\buffer[10][1][0] [3]), .QN());
   DFF_X1 \buffer_reg[10][1][0][2]  (.D(\input_filter[1][0] [2]), .CK(n_56_7), 
      .Q(\buffer[10][1][0] [2]), .QN());
   DFF_X1 \buffer_reg[10][1][0][1]  (.D(\input_filter[1][0] [1]), .CK(n_56_7), 
      .Q(\buffer[10][1][0] [1]), .QN());
   DFF_X1 \buffer_reg[10][1][0][0]  (.D(\input_filter[1][0] [0]), .CK(n_56_7), 
      .Q(\buffer[10][1][0] [0]), .QN());
   DFF_X1 \buffer_reg[11][1][0][15]  (.D(\input_filter[1][0] [15]), .CK(n_56_8), 
      .Q(\buffer[11][1][0] [15]), .QN());
   DFF_X1 \buffer_reg[11][1][0][14]  (.D(\input_filter[1][0] [14]), .CK(n_56_8), 
      .Q(\buffer[11][1][0] [14]), .QN());
   DFF_X1 \buffer_reg[11][1][0][13]  (.D(\input_filter[1][0] [13]), .CK(n_56_8), 
      .Q(\buffer[11][1][0] [13]), .QN());
   DFF_X1 \buffer_reg[11][1][0][12]  (.D(\input_filter[1][0] [12]), .CK(n_56_8), 
      .Q(\buffer[11][1][0] [12]), .QN());
   DFF_X1 \buffer_reg[11][1][0][11]  (.D(\input_filter[1][0] [11]), .CK(n_56_8), 
      .Q(\buffer[11][1][0] [11]), .QN());
   DFF_X1 \buffer_reg[11][1][0][10]  (.D(\input_filter[1][0] [10]), .CK(n_56_8), 
      .Q(\buffer[11][1][0] [10]), .QN());
   DFF_X1 \buffer_reg[11][1][0][9]  (.D(\input_filter[1][0] [9]), .CK(n_56_8), 
      .Q(\buffer[11][1][0] [9]), .QN());
   DFF_X1 \buffer_reg[11][1][0][8]  (.D(\input_filter[1][0] [8]), .CK(n_56_8), 
      .Q(\buffer[11][1][0] [8]), .QN());
   DFF_X1 \buffer_reg[11][1][0][7]  (.D(\input_filter[1][0] [7]), .CK(n_56_8), 
      .Q(\buffer[11][1][0] [7]), .QN());
   DFF_X1 \buffer_reg[11][1][0][6]  (.D(\input_filter[1][0] [6]), .CK(n_56_8), 
      .Q(\buffer[11][1][0] [6]), .QN());
   DFF_X1 \buffer_reg[11][1][0][5]  (.D(\input_filter[1][0] [5]), .CK(n_56_8), 
      .Q(\buffer[11][1][0] [5]), .QN());
   DFF_X1 \buffer_reg[11][1][0][4]  (.D(\input_filter[1][0] [4]), .CK(n_56_8), 
      .Q(\buffer[11][1][0] [4]), .QN());
   DFF_X1 \buffer_reg[11][1][0][3]  (.D(\input_filter[1][0] [3]), .CK(n_56_8), 
      .Q(\buffer[11][1][0] [3]), .QN());
   DFF_X1 \buffer_reg[11][1][0][2]  (.D(\input_filter[1][0] [2]), .CK(n_56_8), 
      .Q(\buffer[11][1][0] [2]), .QN());
   DFF_X1 \buffer_reg[11][1][0][1]  (.D(\input_filter[1][0] [1]), .CK(n_56_8), 
      .Q(\buffer[11][1][0] [1]), .QN());
   DFF_X1 \buffer_reg[11][1][0][0]  (.D(\input_filter[1][0] [0]), .CK(n_56_8), 
      .Q(\buffer[11][1][0] [0]), .QN());
   DFF_X1 \buffer_reg[8][1][2][15]  (.D(\input_filter[1][2] [15]), .CK(n_56_5), 
      .Q(\buffer[8][1][2] [15]), .QN());
   DFF_X1 \buffer_reg[8][1][2][14]  (.D(\input_filter[1][2] [14]), .CK(n_56_5), 
      .Q(\buffer[8][1][2] [14]), .QN());
   DFF_X1 \buffer_reg[8][1][2][13]  (.D(\input_filter[1][2] [13]), .CK(n_56_5), 
      .Q(\buffer[8][1][2] [13]), .QN());
   DFF_X1 \buffer_reg[8][1][2][12]  (.D(\input_filter[1][2] [12]), .CK(n_56_5), 
      .Q(\buffer[8][1][2] [12]), .QN());
   DFF_X1 \buffer_reg[8][1][2][11]  (.D(\input_filter[1][2] [11]), .CK(n_56_5), 
      .Q(\buffer[8][1][2] [11]), .QN());
   DFF_X1 \buffer_reg[8][1][2][10]  (.D(\input_filter[1][2] [10]), .CK(n_56_5), 
      .Q(\buffer[8][1][2] [10]), .QN());
   DFF_X1 \buffer_reg[8][1][2][9]  (.D(\input_filter[1][2] [9]), .CK(n_56_5), 
      .Q(\buffer[8][1][2] [9]), .QN());
   DFF_X1 \buffer_reg[8][1][2][8]  (.D(\input_filter[1][2] [8]), .CK(n_56_5), 
      .Q(\buffer[8][1][2] [8]), .QN());
   DFF_X1 \buffer_reg[8][1][2][7]  (.D(\input_filter[1][2] [7]), .CK(n_56_5), 
      .Q(\buffer[8][1][2] [7]), .QN());
   DFF_X1 \buffer_reg[8][1][2][6]  (.D(\input_filter[1][2] [6]), .CK(n_56_5), 
      .Q(\buffer[8][1][2] [6]), .QN());
   DFF_X1 \buffer_reg[8][1][2][5]  (.D(\input_filter[1][2] [5]), .CK(n_56_5), 
      .Q(\buffer[8][1][2] [5]), .QN());
   DFF_X1 \buffer_reg[8][1][2][4]  (.D(\input_filter[1][2] [4]), .CK(n_56_5), 
      .Q(\buffer[8][1][2] [4]), .QN());
   DFF_X1 \buffer_reg[8][1][2][3]  (.D(\input_filter[1][2] [3]), .CK(n_56_5), 
      .Q(\buffer[8][1][2] [3]), .QN());
   DFF_X1 \buffer_reg[8][1][2][2]  (.D(\input_filter[1][2] [2]), .CK(n_56_5), 
      .Q(\buffer[8][1][2] [2]), .QN());
   DFF_X1 \buffer_reg[8][1][2][1]  (.D(\input_filter[1][2] [1]), .CK(n_56_5), 
      .Q(\buffer[8][1][2] [1]), .QN());
   DFF_X1 \buffer_reg[8][1][2][0]  (.D(\input_filter[1][2] [0]), .CK(n_56_5), 
      .Q(\buffer[8][1][2] [0]), .QN());
   DFF_X1 \buffer_reg[7][1][2][15]  (.D(\input_filter[1][2] [15]), .CK(n_56_4), 
      .Q(\buffer[7][1][2] [15]), .QN());
   DFF_X1 \buffer_reg[7][1][2][14]  (.D(\input_filter[1][2] [14]), .CK(n_56_4), 
      .Q(\buffer[7][1][2] [14]), .QN());
   DFF_X1 \buffer_reg[7][1][2][13]  (.D(\input_filter[1][2] [13]), .CK(n_56_4), 
      .Q(\buffer[7][1][2] [13]), .QN());
   DFF_X1 \buffer_reg[7][1][2][12]  (.D(\input_filter[1][2] [12]), .CK(n_56_4), 
      .Q(\buffer[7][1][2] [12]), .QN());
   DFF_X1 \buffer_reg[7][1][2][11]  (.D(\input_filter[1][2] [11]), .CK(n_56_4), 
      .Q(\buffer[7][1][2] [11]), .QN());
   DFF_X1 \buffer_reg[7][1][2][10]  (.D(\input_filter[1][2] [10]), .CK(n_56_4), 
      .Q(\buffer[7][1][2] [10]), .QN());
   DFF_X1 \buffer_reg[7][1][2][9]  (.D(\input_filter[1][2] [9]), .CK(n_56_4), 
      .Q(\buffer[7][1][2] [9]), .QN());
   DFF_X1 \buffer_reg[7][1][2][8]  (.D(\input_filter[1][2] [8]), .CK(n_56_4), 
      .Q(\buffer[7][1][2] [8]), .QN());
   DFF_X1 \buffer_reg[7][1][2][7]  (.D(\input_filter[1][2] [7]), .CK(n_56_4), 
      .Q(\buffer[7][1][2] [7]), .QN());
   DFF_X1 \buffer_reg[7][1][2][6]  (.D(\input_filter[1][2] [6]), .CK(n_56_4), 
      .Q(\buffer[7][1][2] [6]), .QN());
   DFF_X1 \buffer_reg[7][1][2][5]  (.D(\input_filter[1][2] [5]), .CK(n_56_4), 
      .Q(\buffer[7][1][2] [5]), .QN());
   DFF_X1 \buffer_reg[7][1][2][4]  (.D(\input_filter[1][2] [4]), .CK(n_56_4), 
      .Q(\buffer[7][1][2] [4]), .QN());
   DFF_X1 \buffer_reg[7][1][2][3]  (.D(\input_filter[1][2] [3]), .CK(n_56_4), 
      .Q(\buffer[7][1][2] [3]), .QN());
   DFF_X1 \buffer_reg[7][1][2][2]  (.D(\input_filter[1][2] [2]), .CK(n_56_4), 
      .Q(\buffer[7][1][2] [2]), .QN());
   DFF_X1 \buffer_reg[7][1][2][1]  (.D(\input_filter[1][2] [1]), .CK(n_56_4), 
      .Q(\buffer[7][1][2] [1]), .QN());
   DFF_X1 \buffer_reg[7][1][2][0]  (.D(\input_filter[1][2] [0]), .CK(n_56_4), 
      .Q(\buffer[7][1][2] [0]), .QN());
   DFF_X1 \buffer_reg[6][1][2][15]  (.D(\input_filter[1][2] [15]), .CK(n_56_3), 
      .Q(\buffer[6][1][2] [15]), .QN());
   DFF_X1 \buffer_reg[6][1][2][14]  (.D(\input_filter[1][2] [14]), .CK(n_56_3), 
      .Q(\buffer[6][1][2] [14]), .QN());
   DFF_X1 \buffer_reg[6][1][2][13]  (.D(\input_filter[1][2] [13]), .CK(n_56_3), 
      .Q(\buffer[6][1][2] [13]), .QN());
   DFF_X1 \buffer_reg[6][1][2][12]  (.D(\input_filter[1][2] [12]), .CK(n_56_3), 
      .Q(\buffer[6][1][2] [12]), .QN());
   DFF_X1 \buffer_reg[6][1][2][11]  (.D(\input_filter[1][2] [11]), .CK(n_56_3), 
      .Q(\buffer[6][1][2] [11]), .QN());
   DFF_X1 \buffer_reg[6][1][2][10]  (.D(\input_filter[1][2] [10]), .CK(n_56_3), 
      .Q(\buffer[6][1][2] [10]), .QN());
   DFF_X1 \buffer_reg[6][1][2][9]  (.D(\input_filter[1][2] [9]), .CK(n_56_3), 
      .Q(\buffer[6][1][2] [9]), .QN());
   DFF_X1 \buffer_reg[6][1][2][8]  (.D(\input_filter[1][2] [8]), .CK(n_56_3), 
      .Q(\buffer[6][1][2] [8]), .QN());
   DFF_X1 \buffer_reg[6][1][2][7]  (.D(\input_filter[1][2] [7]), .CK(n_56_3), 
      .Q(\buffer[6][1][2] [7]), .QN());
   DFF_X1 \buffer_reg[6][1][2][6]  (.D(\input_filter[1][2] [6]), .CK(n_56_3), 
      .Q(\buffer[6][1][2] [6]), .QN());
   DFF_X1 \buffer_reg[6][1][2][5]  (.D(\input_filter[1][2] [5]), .CK(n_56_3), 
      .Q(\buffer[6][1][2] [5]), .QN());
   DFF_X1 \buffer_reg[6][1][2][4]  (.D(\input_filter[1][2] [4]), .CK(n_56_3), 
      .Q(\buffer[6][1][2] [4]), .QN());
   DFF_X1 \buffer_reg[6][1][2][3]  (.D(\input_filter[1][2] [3]), .CK(n_56_3), 
      .Q(\buffer[6][1][2] [3]), .QN());
   DFF_X1 \buffer_reg[6][1][2][2]  (.D(\input_filter[1][2] [2]), .CK(n_56_3), 
      .Q(\buffer[6][1][2] [2]), .QN());
   DFF_X1 \buffer_reg[6][1][2][1]  (.D(\input_filter[1][2] [1]), .CK(n_56_3), 
      .Q(\buffer[6][1][2] [1]), .QN());
   DFF_X1 \buffer_reg[6][1][2][0]  (.D(\input_filter[1][2] [0]), .CK(n_56_3), 
      .Q(\buffer[6][1][2] [0]), .QN());
   DFF_X1 \buffer_reg[5][1][2][15]  (.D(\input_filter[1][2] [15]), .CK(n_56_2), 
      .Q(\buffer[5][1][2] [15]), .QN());
   DFF_X1 \buffer_reg[5][1][2][14]  (.D(\input_filter[1][2] [14]), .CK(n_56_2), 
      .Q(\buffer[5][1][2] [14]), .QN());
   DFF_X1 \buffer_reg[5][1][2][13]  (.D(\input_filter[1][2] [13]), .CK(n_56_2), 
      .Q(\buffer[5][1][2] [13]), .QN());
   DFF_X1 \buffer_reg[5][1][2][12]  (.D(\input_filter[1][2] [12]), .CK(n_56_2), 
      .Q(\buffer[5][1][2] [12]), .QN());
   DFF_X1 \buffer_reg[5][1][2][11]  (.D(\input_filter[1][2] [11]), .CK(n_56_2), 
      .Q(\buffer[5][1][2] [11]), .QN());
   DFF_X1 \buffer_reg[5][1][2][10]  (.D(\input_filter[1][2] [10]), .CK(n_56_2), 
      .Q(\buffer[5][1][2] [10]), .QN());
   DFF_X1 \buffer_reg[5][1][2][9]  (.D(\input_filter[1][2] [9]), .CK(n_56_2), 
      .Q(\buffer[5][1][2] [9]), .QN());
   DFF_X1 \buffer_reg[5][1][2][8]  (.D(\input_filter[1][2] [8]), .CK(n_56_2), 
      .Q(\buffer[5][1][2] [8]), .QN());
   DFF_X1 \buffer_reg[5][1][2][7]  (.D(\input_filter[1][2] [7]), .CK(n_56_2), 
      .Q(\buffer[5][1][2] [7]), .QN());
   DFF_X1 \buffer_reg[5][1][2][6]  (.D(\input_filter[1][2] [6]), .CK(n_56_2), 
      .Q(\buffer[5][1][2] [6]), .QN());
   DFF_X1 \buffer_reg[5][1][2][5]  (.D(\input_filter[1][2] [5]), .CK(n_56_2), 
      .Q(\buffer[5][1][2] [5]), .QN());
   DFF_X1 \buffer_reg[5][1][2][4]  (.D(\input_filter[1][2] [4]), .CK(n_56_2), 
      .Q(\buffer[5][1][2] [4]), .QN());
   DFF_X1 \buffer_reg[5][1][2][3]  (.D(\input_filter[1][2] [3]), .CK(n_56_2), 
      .Q(\buffer[5][1][2] [3]), .QN());
   DFF_X1 \buffer_reg[5][1][2][2]  (.D(\input_filter[1][2] [2]), .CK(n_56_2), 
      .Q(\buffer[5][1][2] [2]), .QN());
   DFF_X1 \buffer_reg[5][1][2][1]  (.D(\input_filter[1][2] [1]), .CK(n_56_2), 
      .Q(\buffer[5][1][2] [1]), .QN());
   DFF_X1 \buffer_reg[5][1][2][0]  (.D(\input_filter[1][2] [0]), .CK(n_56_2), 
      .Q(\buffer[5][1][2] [0]), .QN());
   DFF_X1 \buffer_reg[4][1][2][15]  (.D(\input_filter[1][2] [15]), .CK(n_56_1), 
      .Q(\buffer[4][1][2] [15]), .QN());
   DFF_X1 \buffer_reg[4][1][2][14]  (.D(\input_filter[1][2] [14]), .CK(n_56_1), 
      .Q(\buffer[4][1][2] [14]), .QN());
   DFF_X1 \buffer_reg[4][1][2][13]  (.D(\input_filter[1][2] [13]), .CK(n_56_1), 
      .Q(\buffer[4][1][2] [13]), .QN());
   DFF_X1 \buffer_reg[4][1][2][12]  (.D(\input_filter[1][2] [12]), .CK(n_56_1), 
      .Q(\buffer[4][1][2] [12]), .QN());
   DFF_X1 \buffer_reg[4][1][2][11]  (.D(\input_filter[1][2] [11]), .CK(n_56_1), 
      .Q(\buffer[4][1][2] [11]), .QN());
   DFF_X1 \buffer_reg[4][1][2][10]  (.D(\input_filter[1][2] [10]), .CK(n_56_1), 
      .Q(\buffer[4][1][2] [10]), .QN());
   DFF_X1 \buffer_reg[4][1][2][9]  (.D(\input_filter[1][2] [9]), .CK(n_56_1), 
      .Q(\buffer[4][1][2] [9]), .QN());
   DFF_X1 \buffer_reg[4][1][2][8]  (.D(\input_filter[1][2] [8]), .CK(n_56_1), 
      .Q(\buffer[4][1][2] [8]), .QN());
   DFF_X1 \buffer_reg[4][1][2][7]  (.D(\input_filter[1][2] [7]), .CK(n_56_1), 
      .Q(\buffer[4][1][2] [7]), .QN());
   DFF_X1 \buffer_reg[4][1][2][6]  (.D(\input_filter[1][2] [6]), .CK(n_56_1), 
      .Q(\buffer[4][1][2] [6]), .QN());
   DFF_X1 \buffer_reg[4][1][2][5]  (.D(\input_filter[1][2] [5]), .CK(n_56_1), 
      .Q(\buffer[4][1][2] [5]), .QN());
   DFF_X1 \buffer_reg[4][1][2][4]  (.D(\input_filter[1][2] [4]), .CK(n_56_1), 
      .Q(\buffer[4][1][2] [4]), .QN());
   DFF_X1 \buffer_reg[4][1][2][3]  (.D(\input_filter[1][2] [3]), .CK(n_56_1), 
      .Q(\buffer[4][1][2] [3]), .QN());
   DFF_X1 \buffer_reg[4][1][2][2]  (.D(\input_filter[1][2] [2]), .CK(n_56_1), 
      .Q(\buffer[4][1][2] [2]), .QN());
   DFF_X1 \buffer_reg[4][1][2][1]  (.D(\input_filter[1][2] [1]), .CK(n_56_1), 
      .Q(\buffer[4][1][2] [1]), .QN());
   DFF_X1 \buffer_reg[4][1][2][0]  (.D(\input_filter[1][2] [0]), .CK(n_56_1), 
      .Q(\buffer[4][1][2] [0]), .QN());
   DFF_X1 \buffer_reg[3][1][2][15]  (.D(\input_filter[1][2] [15]), .CK(n_56_0), 
      .Q(\buffer[3][1][2] [15]), .QN());
   DFF_X1 \buffer_reg[3][1][2][14]  (.D(\input_filter[1][2] [14]), .CK(n_56_0), 
      .Q(\buffer[3][1][2] [14]), .QN());
   DFF_X1 \buffer_reg[3][1][2][13]  (.D(\input_filter[1][2] [13]), .CK(n_56_0), 
      .Q(\buffer[3][1][2] [13]), .QN());
   DFF_X1 \buffer_reg[3][1][2][12]  (.D(\input_filter[1][2] [12]), .CK(n_56_0), 
      .Q(\buffer[3][1][2] [12]), .QN());
   DFF_X1 \buffer_reg[3][1][2][11]  (.D(\input_filter[1][2] [11]), .CK(n_56_0), 
      .Q(\buffer[3][1][2] [11]), .QN());
   DFF_X1 \buffer_reg[3][1][2][10]  (.D(\input_filter[1][2] [10]), .CK(n_56_0), 
      .Q(\buffer[3][1][2] [10]), .QN());
   DFF_X1 \buffer_reg[3][1][2][9]  (.D(\input_filter[1][2] [9]), .CK(n_56_0), 
      .Q(\buffer[3][1][2] [9]), .QN());
   DFF_X1 \buffer_reg[3][1][2][8]  (.D(\input_filter[1][2] [8]), .CK(n_56_0), 
      .Q(\buffer[3][1][2] [8]), .QN());
   DFF_X1 \buffer_reg[3][1][2][7]  (.D(\input_filter[1][2] [7]), .CK(n_56_0), 
      .Q(\buffer[3][1][2] [7]), .QN());
   DFF_X1 \buffer_reg[3][1][2][6]  (.D(\input_filter[1][2] [6]), .CK(n_56_0), 
      .Q(\buffer[3][1][2] [6]), .QN());
   DFF_X1 \buffer_reg[3][1][2][5]  (.D(\input_filter[1][2] [5]), .CK(n_56_0), 
      .Q(\buffer[3][1][2] [5]), .QN());
   DFF_X1 \buffer_reg[3][1][2][4]  (.D(\input_filter[1][2] [4]), .CK(n_56_0), 
      .Q(\buffer[3][1][2] [4]), .QN());
   DFF_X1 \buffer_reg[3][1][2][3]  (.D(\input_filter[1][2] [3]), .CK(n_56_0), 
      .Q(\buffer[3][1][2] [3]), .QN());
   DFF_X1 \buffer_reg[3][1][2][2]  (.D(\input_filter[1][2] [2]), .CK(n_56_0), 
      .Q(\buffer[3][1][2] [2]), .QN());
   DFF_X1 \buffer_reg[3][1][2][1]  (.D(\input_filter[1][2] [1]), .CK(n_56_0), 
      .Q(\buffer[3][1][2] [1]), .QN());
   DFF_X1 \buffer_reg[3][1][2][0]  (.D(\input_filter[1][2] [0]), .CK(n_56_0), 
      .Q(\buffer[3][1][2] [0]), .QN());
   DFF_X1 \buffer_reg[2][1][2][15]  (.D(\input_filter[1][2] [15]), .CK(n_56_14), 
      .Q(\buffer[2][1][2] [15]), .QN());
   DFF_X1 \buffer_reg[2][1][2][14]  (.D(\input_filter[1][2] [14]), .CK(n_56_14), 
      .Q(\buffer[2][1][2] [14]), .QN());
   DFF_X1 \buffer_reg[2][1][2][13]  (.D(\input_filter[1][2] [13]), .CK(n_56_14), 
      .Q(\buffer[2][1][2] [13]), .QN());
   DFF_X1 \buffer_reg[2][1][2][12]  (.D(\input_filter[1][2] [12]), .CK(n_56_14), 
      .Q(\buffer[2][1][2] [12]), .QN());
   DFF_X1 \buffer_reg[2][1][2][11]  (.D(\input_filter[1][2] [11]), .CK(n_56_14), 
      .Q(\buffer[2][1][2] [11]), .QN());
   DFF_X1 \buffer_reg[2][1][2][10]  (.D(\input_filter[1][2] [10]), .CK(n_56_14), 
      .Q(\buffer[2][1][2] [10]), .QN());
   DFF_X1 \buffer_reg[2][1][2][9]  (.D(\input_filter[1][2] [9]), .CK(n_56_14), 
      .Q(\buffer[2][1][2] [9]), .QN());
   DFF_X1 \buffer_reg[2][1][2][8]  (.D(\input_filter[1][2] [8]), .CK(n_56_14), 
      .Q(\buffer[2][1][2] [8]), .QN());
   DFF_X1 \buffer_reg[2][1][2][7]  (.D(\input_filter[1][2] [7]), .CK(n_56_14), 
      .Q(\buffer[2][1][2] [7]), .QN());
   DFF_X1 \buffer_reg[2][1][2][6]  (.D(\input_filter[1][2] [6]), .CK(n_56_14), 
      .Q(\buffer[2][1][2] [6]), .QN());
   DFF_X1 \buffer_reg[2][1][2][5]  (.D(\input_filter[1][2] [5]), .CK(n_56_14), 
      .Q(\buffer[2][1][2] [5]), .QN());
   DFF_X1 \buffer_reg[2][1][2][4]  (.D(\input_filter[1][2] [4]), .CK(n_56_14), 
      .Q(\buffer[2][1][2] [4]), .QN());
   DFF_X1 \buffer_reg[2][1][2][3]  (.D(\input_filter[1][2] [3]), .CK(n_56_14), 
      .Q(\buffer[2][1][2] [3]), .QN());
   DFF_X1 \buffer_reg[2][1][2][2]  (.D(\input_filter[1][2] [2]), .CK(n_56_14), 
      .Q(\buffer[2][1][2] [2]), .QN());
   DFF_X1 \buffer_reg[2][1][2][1]  (.D(\input_filter[1][2] [1]), .CK(n_56_14), 
      .Q(\buffer[2][1][2] [1]), .QN());
   DFF_X1 \buffer_reg[2][1][2][0]  (.D(\input_filter[1][2] [0]), .CK(n_56_14), 
      .Q(\buffer[2][1][2] [0]), .QN());
   DFF_X1 \buffer_reg[1][1][2][15]  (.D(\input_filter[1][2] [15]), .CK(n_56_13), 
      .Q(\buffer[1][1][2] [15]), .QN());
   DFF_X1 \buffer_reg[1][1][2][14]  (.D(\input_filter[1][2] [14]), .CK(n_56_13), 
      .Q(\buffer[1][1][2] [14]), .QN());
   DFF_X1 \buffer_reg[1][1][2][13]  (.D(\input_filter[1][2] [13]), .CK(n_56_13), 
      .Q(\buffer[1][1][2] [13]), .QN());
   DFF_X1 \buffer_reg[1][1][2][12]  (.D(\input_filter[1][2] [12]), .CK(n_56_13), 
      .Q(\buffer[1][1][2] [12]), .QN());
   DFF_X1 \buffer_reg[1][1][2][11]  (.D(\input_filter[1][2] [11]), .CK(n_56_13), 
      .Q(\buffer[1][1][2] [11]), .QN());
   DFF_X1 \buffer_reg[1][1][2][10]  (.D(\input_filter[1][2] [10]), .CK(n_56_13), 
      .Q(\buffer[1][1][2] [10]), .QN());
   DFF_X1 \buffer_reg[1][1][2][9]  (.D(\input_filter[1][2] [9]), .CK(n_56_13), 
      .Q(\buffer[1][1][2] [9]), .QN());
   DFF_X1 \buffer_reg[1][1][2][8]  (.D(\input_filter[1][2] [8]), .CK(n_56_13), 
      .Q(\buffer[1][1][2] [8]), .QN());
   DFF_X1 \buffer_reg[1][1][2][7]  (.D(\input_filter[1][2] [7]), .CK(n_56_13), 
      .Q(\buffer[1][1][2] [7]), .QN());
   DFF_X1 \buffer_reg[1][1][2][6]  (.D(\input_filter[1][2] [6]), .CK(n_56_13), 
      .Q(\buffer[1][1][2] [6]), .QN());
   DFF_X1 \buffer_reg[1][1][2][5]  (.D(\input_filter[1][2] [5]), .CK(n_56_13), 
      .Q(\buffer[1][1][2] [5]), .QN());
   DFF_X1 \buffer_reg[1][1][2][4]  (.D(\input_filter[1][2] [4]), .CK(n_56_13), 
      .Q(\buffer[1][1][2] [4]), .QN());
   DFF_X1 \buffer_reg[1][1][2][3]  (.D(\input_filter[1][2] [3]), .CK(n_56_13), 
      .Q(\buffer[1][1][2] [3]), .QN());
   DFF_X1 \buffer_reg[1][1][2][2]  (.D(\input_filter[1][2] [2]), .CK(n_56_13), 
      .Q(\buffer[1][1][2] [2]), .QN());
   DFF_X1 \buffer_reg[1][1][2][1]  (.D(\input_filter[1][2] [1]), .CK(n_56_13), 
      .Q(\buffer[1][1][2] [1]), .QN());
   DFF_X1 \buffer_reg[1][1][2][0]  (.D(\input_filter[1][2] [0]), .CK(n_56_13), 
      .Q(\buffer[1][1][2] [0]), .QN());
   DFF_X1 \buffer_reg[12][1][0][15]  (.D(\input_filter[1][0] [15]), .CK(n_56_9), 
      .Q(\buffer[12][1][0] [15]), .QN());
   DFF_X1 \buffer_reg[12][1][0][14]  (.D(\input_filter[1][0] [14]), .CK(n_56_9), 
      .Q(\buffer[12][1][0] [14]), .QN());
   DFF_X1 \buffer_reg[12][1][0][13]  (.D(\input_filter[1][0] [13]), .CK(n_56_9), 
      .Q(\buffer[12][1][0] [13]), .QN());
   DFF_X1 \buffer_reg[12][1][0][12]  (.D(\input_filter[1][0] [12]), .CK(n_56_9), 
      .Q(\buffer[12][1][0] [12]), .QN());
   DFF_X1 \buffer_reg[12][1][0][11]  (.D(\input_filter[1][0] [11]), .CK(n_56_9), 
      .Q(\buffer[12][1][0] [11]), .QN());
   DFF_X1 \buffer_reg[12][1][0][10]  (.D(\input_filter[1][0] [10]), .CK(n_56_9), 
      .Q(\buffer[12][1][0] [10]), .QN());
   DFF_X1 \buffer_reg[12][1][0][9]  (.D(\input_filter[1][0] [9]), .CK(n_56_9), 
      .Q(\buffer[12][1][0] [9]), .QN());
   DFF_X1 \buffer_reg[12][1][0][8]  (.D(\input_filter[1][0] [8]), .CK(n_56_9), 
      .Q(\buffer[12][1][0] [8]), .QN());
   DFF_X1 \buffer_reg[12][1][0][7]  (.D(\input_filter[1][0] [7]), .CK(n_56_9), 
      .Q(\buffer[12][1][0] [7]), .QN());
   DFF_X1 \buffer_reg[12][1][0][6]  (.D(\input_filter[1][0] [6]), .CK(n_56_9), 
      .Q(\buffer[12][1][0] [6]), .QN());
   DFF_X1 \buffer_reg[12][1][0][5]  (.D(\input_filter[1][0] [5]), .CK(n_56_9), 
      .Q(\buffer[12][1][0] [5]), .QN());
   DFF_X1 \buffer_reg[12][1][0][4]  (.D(\input_filter[1][0] [4]), .CK(n_56_9), 
      .Q(\buffer[12][1][0] [4]), .QN());
   DFF_X1 \buffer_reg[12][1][0][3]  (.D(\input_filter[1][0] [3]), .CK(n_56_9), 
      .Q(\buffer[12][1][0] [3]), .QN());
   DFF_X1 \buffer_reg[12][1][0][2]  (.D(\input_filter[1][0] [2]), .CK(n_56_9), 
      .Q(\buffer[12][1][0] [2]), .QN());
   DFF_X1 \buffer_reg[12][1][0][1]  (.D(\input_filter[1][0] [1]), .CK(n_56_9), 
      .Q(\buffer[12][1][0] [1]), .QN());
   DFF_X1 \buffer_reg[12][1][0][0]  (.D(\input_filter[1][0] [0]), .CK(n_56_9), 
      .Q(\buffer[12][1][0] [0]), .QN());
   DFF_X1 \buffer_reg[15][1][1][15]  (.D(\input_filter[1][1] [15]), .CK(n_56_15), 
      .Q(\buffer[15][1][1] [15]), .QN());
   DFF_X1 \buffer_reg[15][1][1][14]  (.D(\input_filter[1][1] [14]), .CK(n_56_15), 
      .Q(\buffer[15][1][1] [14]), .QN());
   DFF_X1 \buffer_reg[15][1][1][13]  (.D(\input_filter[1][1] [13]), .CK(n_56_15), 
      .Q(\buffer[15][1][1] [13]), .QN());
   DFF_X1 \buffer_reg[15][1][1][12]  (.D(\input_filter[1][1] [12]), .CK(n_56_15), 
      .Q(\buffer[15][1][1] [12]), .QN());
   DFF_X1 \buffer_reg[15][1][1][11]  (.D(\input_filter[1][1] [11]), .CK(n_56_15), 
      .Q(\buffer[15][1][1] [11]), .QN());
   DFF_X1 \buffer_reg[15][1][1][10]  (.D(\input_filter[1][1] [10]), .CK(n_56_15), 
      .Q(\buffer[15][1][1] [10]), .QN());
   DFF_X1 \buffer_reg[15][1][1][9]  (.D(\input_filter[1][1] [9]), .CK(n_56_15), 
      .Q(\buffer[15][1][1] [9]), .QN());
   DFF_X1 \buffer_reg[15][1][1][8]  (.D(\input_filter[1][1] [8]), .CK(n_56_15), 
      .Q(\buffer[15][1][1] [8]), .QN());
   DFF_X1 \buffer_reg[15][1][1][7]  (.D(\input_filter[1][1] [7]), .CK(n_56_15), 
      .Q(\buffer[15][1][1] [7]), .QN());
   DFF_X1 \buffer_reg[15][1][1][6]  (.D(\input_filter[1][1] [6]), .CK(n_56_15), 
      .Q(\buffer[15][1][1] [6]), .QN());
   DFF_X1 \buffer_reg[15][1][1][5]  (.D(\input_filter[1][1] [5]), .CK(n_56_15), 
      .Q(\buffer[15][1][1] [5]), .QN());
   DFF_X1 \buffer_reg[15][1][1][4]  (.D(\input_filter[1][1] [4]), .CK(n_56_15), 
      .Q(\buffer[15][1][1] [4]), .QN());
   DFF_X1 \buffer_reg[15][1][1][3]  (.D(\input_filter[1][1] [3]), .CK(n_56_15), 
      .Q(\buffer[15][1][1] [3]), .QN());
   DFF_X1 \buffer_reg[15][1][1][2]  (.D(\input_filter[1][1] [2]), .CK(n_56_15), 
      .Q(\buffer[15][1][1] [2]), .QN());
   DFF_X1 \buffer_reg[15][1][1][1]  (.D(\input_filter[1][1] [1]), .CK(n_56_15), 
      .Q(\buffer[15][1][1] [1]), .QN());
   DFF_X1 \buffer_reg[15][1][1][0]  (.D(\input_filter[1][1] [0]), .CK(n_56_15), 
      .Q(\buffer[15][1][1] [0]), .QN());
   DFF_X1 \buffer_reg[14][1][1][15]  (.D(\input_filter[1][1] [15]), .CK(n_56_11), 
      .Q(\buffer[14][1][1] [15]), .QN());
   DFF_X1 \buffer_reg[14][1][1][14]  (.D(\input_filter[1][1] [14]), .CK(n_56_11), 
      .Q(\buffer[14][1][1] [14]), .QN());
   DFF_X1 \buffer_reg[14][1][1][13]  (.D(\input_filter[1][1] [13]), .CK(n_56_11), 
      .Q(\buffer[14][1][1] [13]), .QN());
   DFF_X1 \buffer_reg[14][1][1][12]  (.D(\input_filter[1][1] [12]), .CK(n_56_11), 
      .Q(\buffer[14][1][1] [12]), .QN());
   DFF_X1 \buffer_reg[14][1][1][11]  (.D(\input_filter[1][1] [11]), .CK(n_56_11), 
      .Q(\buffer[14][1][1] [11]), .QN());
   DFF_X1 \buffer_reg[14][1][1][10]  (.D(\input_filter[1][1] [10]), .CK(n_56_11), 
      .Q(\buffer[14][1][1] [10]), .QN());
   DFF_X1 \buffer_reg[14][1][1][9]  (.D(\input_filter[1][1] [9]), .CK(n_56_11), 
      .Q(\buffer[14][1][1] [9]), .QN());
   DFF_X1 \buffer_reg[14][1][1][8]  (.D(\input_filter[1][1] [8]), .CK(n_56_11), 
      .Q(\buffer[14][1][1] [8]), .QN());
   DFF_X1 \buffer_reg[14][1][1][7]  (.D(\input_filter[1][1] [7]), .CK(n_56_11), 
      .Q(\buffer[14][1][1] [7]), .QN());
   DFF_X1 \buffer_reg[14][1][1][6]  (.D(\input_filter[1][1] [6]), .CK(n_56_11), 
      .Q(\buffer[14][1][1] [6]), .QN());
   DFF_X1 \buffer_reg[14][1][1][5]  (.D(\input_filter[1][1] [5]), .CK(n_56_11), 
      .Q(\buffer[14][1][1] [5]), .QN());
   DFF_X1 \buffer_reg[14][1][1][4]  (.D(\input_filter[1][1] [4]), .CK(n_56_11), 
      .Q(\buffer[14][1][1] [4]), .QN());
   DFF_X1 \buffer_reg[14][1][1][3]  (.D(\input_filter[1][1] [3]), .CK(n_56_11), 
      .Q(\buffer[14][1][1] [3]), .QN());
   DFF_X1 \buffer_reg[14][1][1][2]  (.D(\input_filter[1][1] [2]), .CK(n_56_11), 
      .Q(\buffer[14][1][1] [2]), .QN());
   DFF_X1 \buffer_reg[14][1][1][1]  (.D(\input_filter[1][1] [1]), .CK(n_56_11), 
      .Q(\buffer[14][1][1] [1]), .QN());
   DFF_X1 \buffer_reg[14][1][1][0]  (.D(\input_filter[1][1] [0]), .CK(n_56_11), 
      .Q(\buffer[14][1][1] [0]), .QN());
   DFF_X1 \buffer_reg[13][1][1][15]  (.D(\input_filter[1][1] [15]), .CK(n_56_10), 
      .Q(\buffer[13][1][1] [15]), .QN());
   DFF_X1 \buffer_reg[13][1][1][14]  (.D(\input_filter[1][1] [14]), .CK(n_56_10), 
      .Q(\buffer[13][1][1] [14]), .QN());
   DFF_X1 \buffer_reg[13][1][1][13]  (.D(\input_filter[1][1] [13]), .CK(n_56_10), 
      .Q(\buffer[13][1][1] [13]), .QN());
   DFF_X1 \buffer_reg[13][1][1][12]  (.D(\input_filter[1][1] [12]), .CK(n_56_10), 
      .Q(\buffer[13][1][1] [12]), .QN());
   DFF_X1 \buffer_reg[13][1][1][11]  (.D(\input_filter[1][1] [11]), .CK(n_56_10), 
      .Q(\buffer[13][1][1] [11]), .QN());
   DFF_X1 \buffer_reg[13][1][1][10]  (.D(\input_filter[1][1] [10]), .CK(n_56_10), 
      .Q(\buffer[13][1][1] [10]), .QN());
   DFF_X1 \buffer_reg[13][1][1][9]  (.D(\input_filter[1][1] [9]), .CK(n_56_10), 
      .Q(\buffer[13][1][1] [9]), .QN());
   DFF_X1 \buffer_reg[13][1][1][8]  (.D(\input_filter[1][1] [8]), .CK(n_56_10), 
      .Q(\buffer[13][1][1] [8]), .QN());
   DFF_X1 \buffer_reg[13][1][1][7]  (.D(\input_filter[1][1] [7]), .CK(n_56_10), 
      .Q(\buffer[13][1][1] [7]), .QN());
   DFF_X1 \buffer_reg[13][1][1][6]  (.D(\input_filter[1][1] [6]), .CK(n_56_10), 
      .Q(\buffer[13][1][1] [6]), .QN());
   DFF_X1 \buffer_reg[13][1][1][5]  (.D(\input_filter[1][1] [5]), .CK(n_56_10), 
      .Q(\buffer[13][1][1] [5]), .QN());
   DFF_X1 \buffer_reg[13][1][1][4]  (.D(\input_filter[1][1] [4]), .CK(n_56_10), 
      .Q(\buffer[13][1][1] [4]), .QN());
   DFF_X1 \buffer_reg[13][1][1][3]  (.D(\input_filter[1][1] [3]), .CK(n_56_10), 
      .Q(\buffer[13][1][1] [3]), .QN());
   DFF_X1 \buffer_reg[13][1][1][2]  (.D(\input_filter[1][1] [2]), .CK(n_56_10), 
      .Q(\buffer[13][1][1] [2]), .QN());
   DFF_X1 \buffer_reg[13][1][1][1]  (.D(\input_filter[1][1] [1]), .CK(n_56_10), 
      .Q(\buffer[13][1][1] [1]), .QN());
   DFF_X1 \buffer_reg[13][1][1][0]  (.D(\input_filter[1][1] [0]), .CK(n_56_10), 
      .Q(\buffer[13][1][1] [0]), .QN());
   DFF_X1 \buffer_reg[12][1][1][15]  (.D(\input_filter[1][1] [15]), .CK(n_56_9), 
      .Q(\buffer[12][1][1] [15]), .QN());
   DFF_X1 \buffer_reg[12][1][1][14]  (.D(\input_filter[1][1] [14]), .CK(n_56_9), 
      .Q(\buffer[12][1][1] [14]), .QN());
   DFF_X1 \buffer_reg[12][1][1][13]  (.D(\input_filter[1][1] [13]), .CK(n_56_9), 
      .Q(\buffer[12][1][1] [13]), .QN());
   DFF_X1 \buffer_reg[12][1][1][12]  (.D(\input_filter[1][1] [12]), .CK(n_56_9), 
      .Q(\buffer[12][1][1] [12]), .QN());
   DFF_X1 \buffer_reg[12][1][1][11]  (.D(\input_filter[1][1] [11]), .CK(n_56_9), 
      .Q(\buffer[12][1][1] [11]), .QN());
   DFF_X1 \buffer_reg[12][1][1][10]  (.D(\input_filter[1][1] [10]), .CK(n_56_9), 
      .Q(\buffer[12][1][1] [10]), .QN());
   DFF_X1 \buffer_reg[12][1][1][9]  (.D(\input_filter[1][1] [9]), .CK(n_56_9), 
      .Q(\buffer[12][1][1] [9]), .QN());
   DFF_X1 \buffer_reg[12][1][1][8]  (.D(\input_filter[1][1] [8]), .CK(n_56_9), 
      .Q(\buffer[12][1][1] [8]), .QN());
   DFF_X1 \buffer_reg[12][1][1][7]  (.D(\input_filter[1][1] [7]), .CK(n_56_9), 
      .Q(\buffer[12][1][1] [7]), .QN());
   DFF_X1 \buffer_reg[12][1][1][6]  (.D(\input_filter[1][1] [6]), .CK(n_56_9), 
      .Q(\buffer[12][1][1] [6]), .QN());
   DFF_X1 \buffer_reg[12][1][1][5]  (.D(\input_filter[1][1] [5]), .CK(n_56_9), 
      .Q(\buffer[12][1][1] [5]), .QN());
   DFF_X1 \buffer_reg[12][1][1][4]  (.D(\input_filter[1][1] [4]), .CK(n_56_9), 
      .Q(\buffer[12][1][1] [4]), .QN());
   DFF_X1 \buffer_reg[12][1][1][3]  (.D(\input_filter[1][1] [3]), .CK(n_56_9), 
      .Q(\buffer[12][1][1] [3]), .QN());
   DFF_X1 \buffer_reg[12][1][1][2]  (.D(\input_filter[1][1] [2]), .CK(n_56_9), 
      .Q(\buffer[12][1][1] [2]), .QN());
   DFF_X1 \buffer_reg[12][1][1][1]  (.D(\input_filter[1][1] [1]), .CK(n_56_9), 
      .Q(\buffer[12][1][1] [1]), .QN());
   DFF_X1 \buffer_reg[12][1][1][0]  (.D(\input_filter[1][1] [0]), .CK(n_56_9), 
      .Q(\buffer[12][1][1] [0]), .QN());
   DFF_X1 \buffer_reg[11][1][1][15]  (.D(\input_filter[1][1] [15]), .CK(n_56_8), 
      .Q(\buffer[11][1][1] [15]), .QN());
   DFF_X1 \buffer_reg[11][1][1][14]  (.D(\input_filter[1][1] [14]), .CK(n_56_8), 
      .Q(\buffer[11][1][1] [14]), .QN());
   DFF_X1 \buffer_reg[11][1][1][13]  (.D(\input_filter[1][1] [13]), .CK(n_56_8), 
      .Q(\buffer[11][1][1] [13]), .QN());
   DFF_X1 \buffer_reg[11][1][1][12]  (.D(\input_filter[1][1] [12]), .CK(n_56_8), 
      .Q(\buffer[11][1][1] [12]), .QN());
   DFF_X1 \buffer_reg[11][1][1][11]  (.D(\input_filter[1][1] [11]), .CK(n_56_8), 
      .Q(\buffer[11][1][1] [11]), .QN());
   DFF_X1 \buffer_reg[11][1][1][10]  (.D(\input_filter[1][1] [10]), .CK(n_56_8), 
      .Q(\buffer[11][1][1] [10]), .QN());
   DFF_X1 \buffer_reg[11][1][1][9]  (.D(\input_filter[1][1] [9]), .CK(n_56_8), 
      .Q(\buffer[11][1][1] [9]), .QN());
   DFF_X1 \buffer_reg[11][1][1][8]  (.D(\input_filter[1][1] [8]), .CK(n_56_8), 
      .Q(\buffer[11][1][1] [8]), .QN());
   DFF_X1 \buffer_reg[11][1][1][7]  (.D(\input_filter[1][1] [7]), .CK(n_56_8), 
      .Q(\buffer[11][1][1] [7]), .QN());
   DFF_X1 \buffer_reg[11][1][1][6]  (.D(\input_filter[1][1] [6]), .CK(n_56_8), 
      .Q(\buffer[11][1][1] [6]), .QN());
   DFF_X1 \buffer_reg[11][1][1][5]  (.D(\input_filter[1][1] [5]), .CK(n_56_8), 
      .Q(\buffer[11][1][1] [5]), .QN());
   DFF_X1 \buffer_reg[11][1][1][4]  (.D(\input_filter[1][1] [4]), .CK(n_56_8), 
      .Q(\buffer[11][1][1] [4]), .QN());
   DFF_X1 \buffer_reg[11][1][1][3]  (.D(\input_filter[1][1] [3]), .CK(n_56_8), 
      .Q(\buffer[11][1][1] [3]), .QN());
   DFF_X1 \buffer_reg[11][1][1][2]  (.D(\input_filter[1][1] [2]), .CK(n_56_8), 
      .Q(\buffer[11][1][1] [2]), .QN());
   DFF_X1 \buffer_reg[11][1][1][1]  (.D(\input_filter[1][1] [1]), .CK(n_56_8), 
      .Q(\buffer[11][1][1] [1]), .QN());
   DFF_X1 \buffer_reg[11][1][1][0]  (.D(\input_filter[1][1] [0]), .CK(n_56_8), 
      .Q(\buffer[11][1][1] [0]), .QN());
   DFF_X1 \buffer_reg[10][1][1][15]  (.D(\input_filter[1][1] [15]), .CK(n_56_7), 
      .Q(\buffer[10][1][1] [15]), .QN());
   DFF_X1 \buffer_reg[10][1][1][14]  (.D(\input_filter[1][1] [14]), .CK(n_56_7), 
      .Q(\buffer[10][1][1] [14]), .QN());
   DFF_X1 \buffer_reg[10][1][1][13]  (.D(\input_filter[1][1] [13]), .CK(n_56_7), 
      .Q(\buffer[10][1][1] [13]), .QN());
   DFF_X1 \buffer_reg[10][1][1][12]  (.D(\input_filter[1][1] [12]), .CK(n_56_7), 
      .Q(\buffer[10][1][1] [12]), .QN());
   DFF_X1 \buffer_reg[10][1][1][11]  (.D(\input_filter[1][1] [11]), .CK(n_56_7), 
      .Q(\buffer[10][1][1] [11]), .QN());
   DFF_X1 \buffer_reg[10][1][1][10]  (.D(\input_filter[1][1] [10]), .CK(n_56_7), 
      .Q(\buffer[10][1][1] [10]), .QN());
   DFF_X1 \buffer_reg[10][1][1][9]  (.D(\input_filter[1][1] [9]), .CK(n_56_7), 
      .Q(\buffer[10][1][1] [9]), .QN());
   DFF_X1 \buffer_reg[10][1][1][8]  (.D(\input_filter[1][1] [8]), .CK(n_56_7), 
      .Q(\buffer[10][1][1] [8]), .QN());
   DFF_X1 \buffer_reg[10][1][1][7]  (.D(\input_filter[1][1] [7]), .CK(n_56_7), 
      .Q(\buffer[10][1][1] [7]), .QN());
   DFF_X1 \buffer_reg[10][1][1][6]  (.D(\input_filter[1][1] [6]), .CK(n_56_7), 
      .Q(\buffer[10][1][1] [6]), .QN());
   DFF_X1 \buffer_reg[10][1][1][5]  (.D(\input_filter[1][1] [5]), .CK(n_56_7), 
      .Q(\buffer[10][1][1] [5]), .QN());
   DFF_X1 \buffer_reg[10][1][1][4]  (.D(\input_filter[1][1] [4]), .CK(n_56_7), 
      .Q(\buffer[10][1][1] [4]), .QN());
   DFF_X1 \buffer_reg[10][1][1][3]  (.D(\input_filter[1][1] [3]), .CK(n_56_7), 
      .Q(\buffer[10][1][1] [3]), .QN());
   DFF_X1 \buffer_reg[10][1][1][2]  (.D(\input_filter[1][1] [2]), .CK(n_56_7), 
      .Q(\buffer[10][1][1] [2]), .QN());
   DFF_X1 \buffer_reg[10][1][1][1]  (.D(\input_filter[1][1] [1]), .CK(n_56_7), 
      .Q(\buffer[10][1][1] [1]), .QN());
   DFF_X1 \buffer_reg[10][1][1][0]  (.D(\input_filter[1][1] [0]), .CK(n_56_7), 
      .Q(\buffer[10][1][1] [0]), .QN());
   DFF_X1 \buffer_reg[9][1][1][15]  (.D(\input_filter[1][1] [15]), .CK(n_56_6), 
      .Q(\buffer[9][1][1] [15]), .QN());
   DFF_X1 \buffer_reg[9][1][1][14]  (.D(\input_filter[1][1] [14]), .CK(n_56_6), 
      .Q(\buffer[9][1][1] [14]), .QN());
   DFF_X1 \buffer_reg[9][1][1][13]  (.D(\input_filter[1][1] [13]), .CK(n_56_6), 
      .Q(\buffer[9][1][1] [13]), .QN());
   DFF_X1 \buffer_reg[9][1][1][12]  (.D(\input_filter[1][1] [12]), .CK(n_56_6), 
      .Q(\buffer[9][1][1] [12]), .QN());
   DFF_X1 \buffer_reg[9][1][1][11]  (.D(\input_filter[1][1] [11]), .CK(n_56_6), 
      .Q(\buffer[9][1][1] [11]), .QN());
   DFF_X1 \buffer_reg[9][1][1][10]  (.D(\input_filter[1][1] [10]), .CK(n_56_6), 
      .Q(\buffer[9][1][1] [10]), .QN());
   DFF_X1 \buffer_reg[9][1][1][9]  (.D(\input_filter[1][1] [9]), .CK(n_56_6), 
      .Q(\buffer[9][1][1] [9]), .QN());
   DFF_X1 \buffer_reg[9][1][1][8]  (.D(\input_filter[1][1] [8]), .CK(n_56_6), 
      .Q(\buffer[9][1][1] [8]), .QN());
   DFF_X1 \buffer_reg[9][1][1][7]  (.D(\input_filter[1][1] [7]), .CK(n_56_6), 
      .Q(\buffer[9][1][1] [7]), .QN());
   DFF_X1 \buffer_reg[9][1][1][6]  (.D(\input_filter[1][1] [6]), .CK(n_56_6), 
      .Q(\buffer[9][1][1] [6]), .QN());
   DFF_X1 \buffer_reg[9][1][1][5]  (.D(\input_filter[1][1] [5]), .CK(n_56_6), 
      .Q(\buffer[9][1][1] [5]), .QN());
   DFF_X1 \buffer_reg[9][1][1][4]  (.D(\input_filter[1][1] [4]), .CK(n_56_6), 
      .Q(\buffer[9][1][1] [4]), .QN());
   DFF_X1 \buffer_reg[9][1][1][3]  (.D(\input_filter[1][1] [3]), .CK(n_56_6), 
      .Q(\buffer[9][1][1] [3]), .QN());
   DFF_X1 \buffer_reg[9][1][1][2]  (.D(\input_filter[1][1] [2]), .CK(n_56_6), 
      .Q(\buffer[9][1][1] [2]), .QN());
   DFF_X1 \buffer_reg[9][1][1][1]  (.D(\input_filter[1][1] [1]), .CK(n_56_6), 
      .Q(\buffer[9][1][1] [1]), .QN());
   DFF_X1 \buffer_reg[9][1][1][0]  (.D(\input_filter[1][1] [0]), .CK(n_56_6), 
      .Q(\buffer[9][1][1] [0]), .QN());
   DFF_X1 \buffer_reg[8][1][1][15]  (.D(\input_filter[1][1] [15]), .CK(n_56_5), 
      .Q(\buffer[8][1][1] [15]), .QN());
   DFF_X1 \buffer_reg[8][1][1][14]  (.D(\input_filter[1][1] [14]), .CK(n_56_5), 
      .Q(\buffer[8][1][1] [14]), .QN());
   DFF_X1 \buffer_reg[8][1][1][13]  (.D(\input_filter[1][1] [13]), .CK(n_56_5), 
      .Q(\buffer[8][1][1] [13]), .QN());
   DFF_X1 \buffer_reg[8][1][1][12]  (.D(\input_filter[1][1] [12]), .CK(n_56_5), 
      .Q(\buffer[8][1][1] [12]), .QN());
   DFF_X1 \buffer_reg[8][1][1][11]  (.D(\input_filter[1][1] [11]), .CK(n_56_5), 
      .Q(\buffer[8][1][1] [11]), .QN());
   DFF_X1 \buffer_reg[8][1][1][10]  (.D(\input_filter[1][1] [10]), .CK(n_56_5), 
      .Q(\buffer[8][1][1] [10]), .QN());
   DFF_X1 \buffer_reg[8][1][1][9]  (.D(\input_filter[1][1] [9]), .CK(n_56_5), 
      .Q(\buffer[8][1][1] [9]), .QN());
   DFF_X1 \buffer_reg[8][1][1][8]  (.D(\input_filter[1][1] [8]), .CK(n_56_5), 
      .Q(\buffer[8][1][1] [8]), .QN());
   DFF_X1 \buffer_reg[8][1][1][7]  (.D(\input_filter[1][1] [7]), .CK(n_56_5), 
      .Q(\buffer[8][1][1] [7]), .QN());
   DFF_X1 \buffer_reg[8][1][1][6]  (.D(\input_filter[1][1] [6]), .CK(n_56_5), 
      .Q(\buffer[8][1][1] [6]), .QN());
   DFF_X1 \buffer_reg[8][1][1][5]  (.D(\input_filter[1][1] [5]), .CK(n_56_5), 
      .Q(\buffer[8][1][1] [5]), .QN());
   DFF_X1 \buffer_reg[8][1][1][4]  (.D(\input_filter[1][1] [4]), .CK(n_56_5), 
      .Q(\buffer[8][1][1] [4]), .QN());
   DFF_X1 \buffer_reg[8][1][1][3]  (.D(\input_filter[1][1] [3]), .CK(n_56_5), 
      .Q(\buffer[8][1][1] [3]), .QN());
   DFF_X1 \buffer_reg[8][1][1][2]  (.D(\input_filter[1][1] [2]), .CK(n_56_5), 
      .Q(\buffer[8][1][1] [2]), .QN());
   DFF_X1 \buffer_reg[8][1][1][1]  (.D(\input_filter[1][1] [1]), .CK(n_56_5), 
      .Q(\buffer[8][1][1] [1]), .QN());
   DFF_X1 \buffer_reg[8][1][1][0]  (.D(\input_filter[1][1] [0]), .CK(n_56_5), 
      .Q(\buffer[8][1][1] [0]), .QN());
   DFF_X1 \buffer_reg[7][1][1][15]  (.D(\input_filter[1][1] [15]), .CK(n_56_4), 
      .Q(\buffer[7][1][1] [15]), .QN());
   DFF_X1 \buffer_reg[7][1][1][14]  (.D(\input_filter[1][1] [14]), .CK(n_56_4), 
      .Q(\buffer[7][1][1] [14]), .QN());
   DFF_X1 \buffer_reg[7][1][1][13]  (.D(\input_filter[1][1] [13]), .CK(n_56_4), 
      .Q(\buffer[7][1][1] [13]), .QN());
   DFF_X1 \buffer_reg[7][1][1][12]  (.D(\input_filter[1][1] [12]), .CK(n_56_4), 
      .Q(\buffer[7][1][1] [12]), .QN());
   DFF_X1 \buffer_reg[7][1][1][11]  (.D(\input_filter[1][1] [11]), .CK(n_56_4), 
      .Q(\buffer[7][1][1] [11]), .QN());
   DFF_X1 \buffer_reg[7][1][1][10]  (.D(\input_filter[1][1] [10]), .CK(n_56_4), 
      .Q(\buffer[7][1][1] [10]), .QN());
   DFF_X1 \buffer_reg[7][1][1][9]  (.D(\input_filter[1][1] [9]), .CK(n_56_4), 
      .Q(\buffer[7][1][1] [9]), .QN());
   DFF_X1 \buffer_reg[7][1][1][8]  (.D(\input_filter[1][1] [8]), .CK(n_56_4), 
      .Q(\buffer[7][1][1] [8]), .QN());
   DFF_X1 \buffer_reg[7][1][1][7]  (.D(\input_filter[1][1] [7]), .CK(n_56_4), 
      .Q(\buffer[7][1][1] [7]), .QN());
   DFF_X1 \buffer_reg[7][1][1][6]  (.D(\input_filter[1][1] [6]), .CK(n_56_4), 
      .Q(\buffer[7][1][1] [6]), .QN());
   DFF_X1 \buffer_reg[7][1][1][5]  (.D(\input_filter[1][1] [5]), .CK(n_56_4), 
      .Q(\buffer[7][1][1] [5]), .QN());
   DFF_X1 \buffer_reg[7][1][1][4]  (.D(\input_filter[1][1] [4]), .CK(n_56_4), 
      .Q(\buffer[7][1][1] [4]), .QN());
   DFF_X1 \buffer_reg[7][1][1][3]  (.D(\input_filter[1][1] [3]), .CK(n_56_4), 
      .Q(\buffer[7][1][1] [3]), .QN());
   DFF_X1 \buffer_reg[7][1][1][2]  (.D(\input_filter[1][1] [2]), .CK(n_56_4), 
      .Q(\buffer[7][1][1] [2]), .QN());
   DFF_X1 \buffer_reg[7][1][1][1]  (.D(\input_filter[1][1] [1]), .CK(n_56_4), 
      .Q(\buffer[7][1][1] [1]), .QN());
   DFF_X1 \buffer_reg[7][1][1][0]  (.D(\input_filter[1][1] [0]), .CK(n_56_4), 
      .Q(\buffer[7][1][1] [0]), .QN());
   DFF_X1 \buffer_reg[6][1][1][15]  (.D(\input_filter[1][1] [15]), .CK(n_56_3), 
      .Q(\buffer[6][1][1] [15]), .QN());
   DFF_X1 \buffer_reg[6][1][1][14]  (.D(\input_filter[1][1] [14]), .CK(n_56_3), 
      .Q(\buffer[6][1][1] [14]), .QN());
   DFF_X1 \buffer_reg[6][1][1][13]  (.D(\input_filter[1][1] [13]), .CK(n_56_3), 
      .Q(\buffer[6][1][1] [13]), .QN());
   DFF_X1 \buffer_reg[6][1][1][12]  (.D(\input_filter[1][1] [12]), .CK(n_56_3), 
      .Q(\buffer[6][1][1] [12]), .QN());
   DFF_X1 \buffer_reg[6][1][1][11]  (.D(\input_filter[1][1] [11]), .CK(n_56_3), 
      .Q(\buffer[6][1][1] [11]), .QN());
   DFF_X1 \buffer_reg[6][1][1][10]  (.D(\input_filter[1][1] [10]), .CK(n_56_3), 
      .Q(\buffer[6][1][1] [10]), .QN());
   DFF_X1 \buffer_reg[6][1][1][9]  (.D(\input_filter[1][1] [9]), .CK(n_56_3), 
      .Q(\buffer[6][1][1] [9]), .QN());
   DFF_X1 \buffer_reg[6][1][1][8]  (.D(\input_filter[1][1] [8]), .CK(n_56_3), 
      .Q(\buffer[6][1][1] [8]), .QN());
   DFF_X1 \buffer_reg[6][1][1][7]  (.D(\input_filter[1][1] [7]), .CK(n_56_3), 
      .Q(\buffer[6][1][1] [7]), .QN());
   DFF_X1 \buffer_reg[6][1][1][6]  (.D(\input_filter[1][1] [6]), .CK(n_56_3), 
      .Q(\buffer[6][1][1] [6]), .QN());
   DFF_X1 \buffer_reg[6][1][1][5]  (.D(\input_filter[1][1] [5]), .CK(n_56_3), 
      .Q(\buffer[6][1][1] [5]), .QN());
   DFF_X1 \buffer_reg[6][1][1][4]  (.D(\input_filter[1][1] [4]), .CK(n_56_3), 
      .Q(\buffer[6][1][1] [4]), .QN());
   DFF_X1 \buffer_reg[6][1][1][3]  (.D(\input_filter[1][1] [3]), .CK(n_56_3), 
      .Q(\buffer[6][1][1] [3]), .QN());
   DFF_X1 \buffer_reg[6][1][1][2]  (.D(\input_filter[1][1] [2]), .CK(n_56_3), 
      .Q(\buffer[6][1][1] [2]), .QN());
   DFF_X1 \buffer_reg[6][1][1][1]  (.D(\input_filter[1][1] [1]), .CK(n_56_3), 
      .Q(\buffer[6][1][1] [1]), .QN());
   DFF_X1 \buffer_reg[6][1][1][0]  (.D(\input_filter[1][1] [0]), .CK(n_56_3), 
      .Q(\buffer[6][1][1] [0]), .QN());
   DFF_X1 \buffer_reg[5][1][1][15]  (.D(\input_filter[1][1] [15]), .CK(n_56_2), 
      .Q(\buffer[5][1][1] [15]), .QN());
   DFF_X1 \buffer_reg[5][1][1][14]  (.D(\input_filter[1][1] [14]), .CK(n_56_2), 
      .Q(\buffer[5][1][1] [14]), .QN());
   DFF_X1 \buffer_reg[5][1][1][13]  (.D(\input_filter[1][1] [13]), .CK(n_56_2), 
      .Q(\buffer[5][1][1] [13]), .QN());
   DFF_X1 \buffer_reg[5][1][1][12]  (.D(\input_filter[1][1] [12]), .CK(n_56_2), 
      .Q(\buffer[5][1][1] [12]), .QN());
   DFF_X1 \buffer_reg[5][1][1][11]  (.D(\input_filter[1][1] [11]), .CK(n_56_2), 
      .Q(\buffer[5][1][1] [11]), .QN());
   DFF_X1 \buffer_reg[5][1][1][10]  (.D(\input_filter[1][1] [10]), .CK(n_56_2), 
      .Q(\buffer[5][1][1] [10]), .QN());
   DFF_X1 \buffer_reg[5][1][1][9]  (.D(\input_filter[1][1] [9]), .CK(n_56_2), 
      .Q(\buffer[5][1][1] [9]), .QN());
   DFF_X1 \buffer_reg[5][1][1][8]  (.D(\input_filter[1][1] [8]), .CK(n_56_2), 
      .Q(\buffer[5][1][1] [8]), .QN());
   DFF_X1 \buffer_reg[5][1][1][7]  (.D(\input_filter[1][1] [7]), .CK(n_56_2), 
      .Q(\buffer[5][1][1] [7]), .QN());
   DFF_X1 \buffer_reg[5][1][1][6]  (.D(\input_filter[1][1] [6]), .CK(n_56_2), 
      .Q(\buffer[5][1][1] [6]), .QN());
   DFF_X1 \buffer_reg[5][1][1][5]  (.D(\input_filter[1][1] [5]), .CK(n_56_2), 
      .Q(\buffer[5][1][1] [5]), .QN());
   DFF_X1 \buffer_reg[5][1][1][4]  (.D(\input_filter[1][1] [4]), .CK(n_56_2), 
      .Q(\buffer[5][1][1] [4]), .QN());
   DFF_X1 \buffer_reg[5][1][1][3]  (.D(\input_filter[1][1] [3]), .CK(n_56_2), 
      .Q(\buffer[5][1][1] [3]), .QN());
   DFF_X1 \buffer_reg[5][1][1][2]  (.D(\input_filter[1][1] [2]), .CK(n_56_2), 
      .Q(\buffer[5][1][1] [2]), .QN());
   DFF_X1 \buffer_reg[5][1][1][1]  (.D(\input_filter[1][1] [1]), .CK(n_56_2), 
      .Q(\buffer[5][1][1] [1]), .QN());
   DFF_X1 \buffer_reg[5][1][1][0]  (.D(\input_filter[1][1] [0]), .CK(n_56_2), 
      .Q(\buffer[5][1][1] [0]), .QN());
   DFF_X1 \buffer_reg[4][1][1][15]  (.D(\input_filter[1][1] [15]), .CK(n_56_1), 
      .Q(\buffer[4][1][1] [15]), .QN());
   DFF_X1 \buffer_reg[4][1][1][14]  (.D(\input_filter[1][1] [14]), .CK(n_56_1), 
      .Q(\buffer[4][1][1] [14]), .QN());
   DFF_X1 \buffer_reg[4][1][1][13]  (.D(\input_filter[1][1] [13]), .CK(n_56_1), 
      .Q(\buffer[4][1][1] [13]), .QN());
   DFF_X1 \buffer_reg[4][1][1][12]  (.D(\input_filter[1][1] [12]), .CK(n_56_1), 
      .Q(\buffer[4][1][1] [12]), .QN());
   DFF_X1 \buffer_reg[4][1][1][11]  (.D(\input_filter[1][1] [11]), .CK(n_56_1), 
      .Q(\buffer[4][1][1] [11]), .QN());
   DFF_X1 \buffer_reg[4][1][1][10]  (.D(\input_filter[1][1] [10]), .CK(n_56_1), 
      .Q(\buffer[4][1][1] [10]), .QN());
   DFF_X1 \buffer_reg[4][1][1][9]  (.D(\input_filter[1][1] [9]), .CK(n_56_1), 
      .Q(\buffer[4][1][1] [9]), .QN());
   DFF_X1 \buffer_reg[4][1][1][8]  (.D(\input_filter[1][1] [8]), .CK(n_56_1), 
      .Q(\buffer[4][1][1] [8]), .QN());
   DFF_X1 \buffer_reg[4][1][1][7]  (.D(\input_filter[1][1] [7]), .CK(n_56_1), 
      .Q(\buffer[4][1][1] [7]), .QN());
   DFF_X1 \buffer_reg[4][1][1][6]  (.D(\input_filter[1][1] [6]), .CK(n_56_1), 
      .Q(\buffer[4][1][1] [6]), .QN());
   DFF_X1 \buffer_reg[4][1][1][5]  (.D(\input_filter[1][1] [5]), .CK(n_56_1), 
      .Q(\buffer[4][1][1] [5]), .QN());
   DFF_X1 \buffer_reg[4][1][1][4]  (.D(\input_filter[1][1] [4]), .CK(n_56_1), 
      .Q(\buffer[4][1][1] [4]), .QN());
   DFF_X1 \buffer_reg[4][1][1][3]  (.D(\input_filter[1][1] [3]), .CK(n_56_1), 
      .Q(\buffer[4][1][1] [3]), .QN());
   DFF_X1 \buffer_reg[4][1][1][2]  (.D(\input_filter[1][1] [2]), .CK(n_56_1), 
      .Q(\buffer[4][1][1] [2]), .QN());
   DFF_X1 \buffer_reg[4][1][1][1]  (.D(\input_filter[1][1] [1]), .CK(n_56_1), 
      .Q(\buffer[4][1][1] [1]), .QN());
   DFF_X1 \buffer_reg[4][1][1][0]  (.D(\input_filter[1][1] [0]), .CK(n_56_1), 
      .Q(\buffer[4][1][1] [0]), .QN());
   DFF_X1 \buffer_reg[3][1][1][15]  (.D(\input_filter[1][1] [15]), .CK(n_56_0), 
      .Q(\buffer[3][1][1] [15]), .QN());
   DFF_X1 \buffer_reg[3][1][1][14]  (.D(\input_filter[1][1] [14]), .CK(n_56_0), 
      .Q(\buffer[3][1][1] [14]), .QN());
   DFF_X1 \buffer_reg[3][1][1][13]  (.D(\input_filter[1][1] [13]), .CK(n_56_0), 
      .Q(\buffer[3][1][1] [13]), .QN());
   DFF_X1 \buffer_reg[3][1][1][12]  (.D(\input_filter[1][1] [12]), .CK(n_56_0), 
      .Q(\buffer[3][1][1] [12]), .QN());
   DFF_X1 \buffer_reg[3][1][1][11]  (.D(\input_filter[1][1] [11]), .CK(n_56_0), 
      .Q(\buffer[3][1][1] [11]), .QN());
   DFF_X1 \buffer_reg[3][1][1][10]  (.D(\input_filter[1][1] [10]), .CK(n_56_0), 
      .Q(\buffer[3][1][1] [10]), .QN());
   DFF_X1 \buffer_reg[3][1][1][9]  (.D(\input_filter[1][1] [9]), .CK(n_56_0), 
      .Q(\buffer[3][1][1] [9]), .QN());
   DFF_X1 \buffer_reg[3][1][1][8]  (.D(\input_filter[1][1] [8]), .CK(n_56_0), 
      .Q(\buffer[3][1][1] [8]), .QN());
   DFF_X1 \buffer_reg[3][1][1][7]  (.D(\input_filter[1][1] [7]), .CK(n_56_0), 
      .Q(\buffer[3][1][1] [7]), .QN());
   DFF_X1 \buffer_reg[3][1][1][6]  (.D(\input_filter[1][1] [6]), .CK(n_56_0), 
      .Q(\buffer[3][1][1] [6]), .QN());
   DFF_X1 \buffer_reg[3][1][1][5]  (.D(\input_filter[1][1] [5]), .CK(n_56_0), 
      .Q(\buffer[3][1][1] [5]), .QN());
   DFF_X1 \buffer_reg[3][1][1][4]  (.D(\input_filter[1][1] [4]), .CK(n_56_0), 
      .Q(\buffer[3][1][1] [4]), .QN());
   DFF_X1 \buffer_reg[3][1][1][3]  (.D(\input_filter[1][1] [3]), .CK(n_56_0), 
      .Q(\buffer[3][1][1] [3]), .QN());
   DFF_X1 \buffer_reg[3][1][1][2]  (.D(\input_filter[1][1] [2]), .CK(n_56_0), 
      .Q(\buffer[3][1][1] [2]), .QN());
   DFF_X1 \buffer_reg[3][1][1][1]  (.D(\input_filter[1][1] [1]), .CK(n_56_0), 
      .Q(\buffer[3][1][1] [1]), .QN());
   DFF_X1 \buffer_reg[3][1][1][0]  (.D(\input_filter[1][1] [0]), .CK(n_56_0), 
      .Q(\buffer[3][1][1] [0]), .QN());
   DFF_X1 \buffer_reg[2][1][1][15]  (.D(\input_filter[1][1] [15]), .CK(n_56_14), 
      .Q(\buffer[2][1][1] [15]), .QN());
   DFF_X1 \buffer_reg[2][1][1][14]  (.D(\input_filter[1][1] [14]), .CK(n_56_14), 
      .Q(\buffer[2][1][1] [14]), .QN());
   DFF_X1 \buffer_reg[2][1][1][13]  (.D(\input_filter[1][1] [13]), .CK(n_56_14), 
      .Q(\buffer[2][1][1] [13]), .QN());
   DFF_X1 \buffer_reg[2][1][1][12]  (.D(\input_filter[1][1] [12]), .CK(n_56_14), 
      .Q(\buffer[2][1][1] [12]), .QN());
   DFF_X1 \buffer_reg[2][1][1][11]  (.D(\input_filter[1][1] [11]), .CK(n_56_14), 
      .Q(\buffer[2][1][1] [11]), .QN());
   DFF_X1 \buffer_reg[2][1][1][10]  (.D(\input_filter[1][1] [10]), .CK(n_56_14), 
      .Q(\buffer[2][1][1] [10]), .QN());
   DFF_X1 \buffer_reg[2][1][1][9]  (.D(\input_filter[1][1] [9]), .CK(n_56_14), 
      .Q(\buffer[2][1][1] [9]), .QN());
   DFF_X1 \buffer_reg[2][1][1][8]  (.D(\input_filter[1][1] [8]), .CK(n_56_14), 
      .Q(\buffer[2][1][1] [8]), .QN());
   DFF_X1 \buffer_reg[2][1][1][7]  (.D(\input_filter[1][1] [7]), .CK(n_56_14), 
      .Q(\buffer[2][1][1] [7]), .QN());
   DFF_X1 \buffer_reg[2][1][1][6]  (.D(\input_filter[1][1] [6]), .CK(n_56_14), 
      .Q(\buffer[2][1][1] [6]), .QN());
   DFF_X1 \buffer_reg[2][1][1][5]  (.D(\input_filter[1][1] [5]), .CK(n_56_14), 
      .Q(\buffer[2][1][1] [5]), .QN());
   DFF_X1 \buffer_reg[2][1][1][4]  (.D(\input_filter[1][1] [4]), .CK(n_56_14), 
      .Q(\buffer[2][1][1] [4]), .QN());
   DFF_X1 \buffer_reg[2][1][1][3]  (.D(\input_filter[1][1] [3]), .CK(n_56_14), 
      .Q(\buffer[2][1][1] [3]), .QN());
   DFF_X1 \buffer_reg[2][1][1][2]  (.D(\input_filter[1][1] [2]), .CK(n_56_14), 
      .Q(\buffer[2][1][1] [2]), .QN());
   DFF_X1 \buffer_reg[2][1][1][1]  (.D(\input_filter[1][1] [1]), .CK(n_56_14), 
      .Q(\buffer[2][1][1] [1]), .QN());
   DFF_X1 \buffer_reg[2][1][1][0]  (.D(\input_filter[1][1] [0]), .CK(n_56_14), 
      .Q(\buffer[2][1][1] [0]), .QN());
   DFF_X1 \buffer_reg[1][1][1][15]  (.D(\input_filter[1][1] [15]), .CK(n_56_13), 
      .Q(\buffer[1][1][1] [15]), .QN());
   DFF_X1 \buffer_reg[1][1][1][14]  (.D(\input_filter[1][1] [14]), .CK(n_56_13), 
      .Q(\buffer[1][1][1] [14]), .QN());
   DFF_X1 \buffer_reg[1][1][1][13]  (.D(\input_filter[1][1] [13]), .CK(n_56_13), 
      .Q(\buffer[1][1][1] [13]), .QN());
   DFF_X1 \buffer_reg[1][1][1][12]  (.D(\input_filter[1][1] [12]), .CK(n_56_13), 
      .Q(\buffer[1][1][1] [12]), .QN());
   DFF_X1 \buffer_reg[1][1][1][11]  (.D(\input_filter[1][1] [11]), .CK(n_56_13), 
      .Q(\buffer[1][1][1] [11]), .QN());
   DFF_X1 \buffer_reg[1][1][1][10]  (.D(\input_filter[1][1] [10]), .CK(n_56_13), 
      .Q(\buffer[1][1][1] [10]), .QN());
   DFF_X1 \buffer_reg[1][1][1][9]  (.D(\input_filter[1][1] [9]), .CK(n_56_13), 
      .Q(\buffer[1][1][1] [9]), .QN());
   DFF_X1 \buffer_reg[1][1][1][8]  (.D(\input_filter[1][1] [8]), .CK(n_56_13), 
      .Q(\buffer[1][1][1] [8]), .QN());
   DFF_X1 \buffer_reg[1][1][1][7]  (.D(\input_filter[1][1] [7]), .CK(n_56_13), 
      .Q(\buffer[1][1][1] [7]), .QN());
   DFF_X1 \buffer_reg[1][1][1][6]  (.D(\input_filter[1][1] [6]), .CK(n_56_13), 
      .Q(\buffer[1][1][1] [6]), .QN());
   DFF_X1 \buffer_reg[1][1][1][5]  (.D(\input_filter[1][1] [5]), .CK(n_56_13), 
      .Q(\buffer[1][1][1] [5]), .QN());
   DFF_X1 \buffer_reg[1][1][1][4]  (.D(\input_filter[1][1] [4]), .CK(n_56_13), 
      .Q(\buffer[1][1][1] [4]), .QN());
   DFF_X1 \buffer_reg[1][1][1][3]  (.D(\input_filter[1][1] [3]), .CK(n_56_13), 
      .Q(\buffer[1][1][1] [3]), .QN());
   DFF_X1 \buffer_reg[1][1][1][2]  (.D(\input_filter[1][1] [2]), .CK(n_56_13), 
      .Q(\buffer[1][1][1] [2]), .QN());
   DFF_X1 \buffer_reg[1][1][1][1]  (.D(\input_filter[1][1] [1]), .CK(n_56_13), 
      .Q(\buffer[1][1][1] [1]), .QN());
   DFF_X1 \buffer_reg[1][1][1][0]  (.D(\input_filter[1][1] [0]), .CK(n_56_13), 
      .Q(\buffer[1][1][1] [0]), .QN());
   DFF_X1 \buffer_reg[0][1][1][15]  (.D(\input_filter[1][1] [15]), .CK(n_56_12), 
      .Q(\buffer[0][1][1] [15]), .QN());
   DFF_X1 \buffer_reg[0][1][1][14]  (.D(\input_filter[1][1] [14]), .CK(n_56_12), 
      .Q(\buffer[0][1][1] [14]), .QN());
   DFF_X1 \buffer_reg[0][1][1][13]  (.D(\input_filter[1][1] [13]), .CK(n_56_12), 
      .Q(\buffer[0][1][1] [13]), .QN());
   DFF_X1 \buffer_reg[0][1][1][12]  (.D(\input_filter[1][1] [12]), .CK(n_56_12), 
      .Q(\buffer[0][1][1] [12]), .QN());
   DFF_X1 \buffer_reg[0][1][1][11]  (.D(\input_filter[1][1] [11]), .CK(n_56_12), 
      .Q(\buffer[0][1][1] [11]), .QN());
   DFF_X1 \buffer_reg[0][1][1][10]  (.D(\input_filter[1][1] [10]), .CK(n_56_12), 
      .Q(\buffer[0][1][1] [10]), .QN());
   DFF_X1 \buffer_reg[0][1][1][9]  (.D(\input_filter[1][1] [9]), .CK(n_56_12), 
      .Q(\buffer[0][1][1] [9]), .QN());
   DFF_X1 \buffer_reg[0][1][1][8]  (.D(\input_filter[1][1] [8]), .CK(n_56_12), 
      .Q(\buffer[0][1][1] [8]), .QN());
   DFF_X1 \buffer_reg[0][1][1][7]  (.D(\input_filter[1][1] [7]), .CK(n_56_12), 
      .Q(\buffer[0][1][1] [7]), .QN());
   DFF_X1 \buffer_reg[0][1][1][6]  (.D(\input_filter[1][1] [6]), .CK(n_56_12), 
      .Q(\buffer[0][1][1] [6]), .QN());
   DFF_X1 \buffer_reg[0][1][1][5]  (.D(\input_filter[1][1] [5]), .CK(n_56_12), 
      .Q(\buffer[0][1][1] [5]), .QN());
   DFF_X1 \buffer_reg[0][1][1][4]  (.D(\input_filter[1][1] [4]), .CK(n_56_12), 
      .Q(\buffer[0][1][1] [4]), .QN());
   DFF_X1 \buffer_reg[0][1][1][3]  (.D(\input_filter[1][1] [3]), .CK(n_56_12), 
      .Q(\buffer[0][1][1] [3]), .QN());
   DFF_X1 \buffer_reg[0][1][1][2]  (.D(\input_filter[1][1] [2]), .CK(n_56_12), 
      .Q(\buffer[0][1][1] [2]), .QN());
   DFF_X1 \buffer_reg[0][1][1][1]  (.D(\input_filter[1][1] [1]), .CK(n_56_12), 
      .Q(\buffer[0][1][1] [1]), .QN());
   DFF_X1 \buffer_reg[0][1][1][0]  (.D(\input_filter[1][1] [0]), .CK(n_56_12), 
      .Q(\buffer[0][1][1] [0]), .QN());
   DFF_X1 \buffer_reg[15][1][0][15]  (.D(\input_filter[1][0] [15]), .CK(n_56_15), 
      .Q(\buffer[15][1][0] [15]), .QN());
   DFF_X1 \buffer_reg[15][1][0][14]  (.D(\input_filter[1][0] [14]), .CK(n_56_15), 
      .Q(\buffer[15][1][0] [14]), .QN());
   DFF_X1 \buffer_reg[15][1][0][13]  (.D(\input_filter[1][0] [13]), .CK(n_56_15), 
      .Q(\buffer[15][1][0] [13]), .QN());
   DFF_X1 \buffer_reg[15][1][0][12]  (.D(\input_filter[1][0] [12]), .CK(n_56_15), 
      .Q(\buffer[15][1][0] [12]), .QN());
   DFF_X1 \buffer_reg[15][1][0][11]  (.D(\input_filter[1][0] [11]), .CK(n_56_15), 
      .Q(\buffer[15][1][0] [11]), .QN());
   DFF_X1 \buffer_reg[15][1][0][10]  (.D(\input_filter[1][0] [10]), .CK(n_56_15), 
      .Q(\buffer[15][1][0] [10]), .QN());
   DFF_X1 \buffer_reg[15][1][0][9]  (.D(\input_filter[1][0] [9]), .CK(n_56_15), 
      .Q(\buffer[15][1][0] [9]), .QN());
   DFF_X1 \buffer_reg[15][1][0][8]  (.D(\input_filter[1][0] [8]), .CK(n_56_15), 
      .Q(\buffer[15][1][0] [8]), .QN());
   DFF_X1 \buffer_reg[15][1][0][7]  (.D(\input_filter[1][0] [7]), .CK(n_56_15), 
      .Q(\buffer[15][1][0] [7]), .QN());
   DFF_X1 \buffer_reg[15][1][0][6]  (.D(\input_filter[1][0] [6]), .CK(n_56_15), 
      .Q(\buffer[15][1][0] [6]), .QN());
   DFF_X1 \buffer_reg[15][1][0][5]  (.D(\input_filter[1][0] [5]), .CK(n_56_15), 
      .Q(\buffer[15][1][0] [5]), .QN());
   DFF_X1 \buffer_reg[15][1][0][4]  (.D(\input_filter[1][0] [4]), .CK(n_56_15), 
      .Q(\buffer[15][1][0] [4]), .QN());
   DFF_X1 \buffer_reg[15][1][0][3]  (.D(\input_filter[1][0] [3]), .CK(n_56_15), 
      .Q(\buffer[15][1][0] [3]), .QN());
   DFF_X1 \buffer_reg[15][1][0][2]  (.D(\input_filter[1][0] [2]), .CK(n_56_15), 
      .Q(\buffer[15][1][0] [2]), .QN());
   DFF_X1 \buffer_reg[15][1][0][1]  (.D(\input_filter[1][0] [1]), .CK(n_56_15), 
      .Q(\buffer[15][1][0] [1]), .QN());
   DFF_X1 \buffer_reg[15][1][0][0]  (.D(\input_filter[1][0] [0]), .CK(n_56_15), 
      .Q(\buffer[15][1][0] [0]), .QN());
   DFF_X1 \buffer_reg[14][1][0][15]  (.D(\input_filter[1][0] [15]), .CK(n_56_11), 
      .Q(\buffer[14][1][0] [15]), .QN());
   DFF_X1 \buffer_reg[14][1][0][14]  (.D(\input_filter[1][0] [14]), .CK(n_56_11), 
      .Q(\buffer[14][1][0] [14]), .QN());
   DFF_X1 \buffer_reg[14][1][0][13]  (.D(\input_filter[1][0] [13]), .CK(n_56_11), 
      .Q(\buffer[14][1][0] [13]), .QN());
   DFF_X1 \buffer_reg[14][1][0][12]  (.D(\input_filter[1][0] [12]), .CK(n_56_11), 
      .Q(\buffer[14][1][0] [12]), .QN());
   DFF_X1 \buffer_reg[14][1][0][11]  (.D(\input_filter[1][0] [11]), .CK(n_56_11), 
      .Q(\buffer[14][1][0] [11]), .QN());
   DFF_X1 \buffer_reg[14][1][0][10]  (.D(\input_filter[1][0] [10]), .CK(n_56_11), 
      .Q(\buffer[14][1][0] [10]), .QN());
   DFF_X1 \buffer_reg[14][1][0][9]  (.D(\input_filter[1][0] [9]), .CK(n_56_11), 
      .Q(\buffer[14][1][0] [9]), .QN());
   DFF_X1 \buffer_reg[14][1][0][8]  (.D(\input_filter[1][0] [8]), .CK(n_56_11), 
      .Q(\buffer[14][1][0] [8]), .QN());
   DFF_X1 \buffer_reg[14][1][0][7]  (.D(\input_filter[1][0] [7]), .CK(n_56_11), 
      .Q(\buffer[14][1][0] [7]), .QN());
   DFF_X1 \buffer_reg[14][1][0][6]  (.D(\input_filter[1][0] [6]), .CK(n_56_11), 
      .Q(\buffer[14][1][0] [6]), .QN());
   DFF_X1 \buffer_reg[14][1][0][5]  (.D(\input_filter[1][0] [5]), .CK(n_56_11), 
      .Q(\buffer[14][1][0] [5]), .QN());
   DFF_X1 \buffer_reg[14][1][0][4]  (.D(\input_filter[1][0] [4]), .CK(n_56_11), 
      .Q(\buffer[14][1][0] [4]), .QN());
   DFF_X1 \buffer_reg[14][1][0][3]  (.D(\input_filter[1][0] [3]), .CK(n_56_11), 
      .Q(\buffer[14][1][0] [3]), .QN());
   DFF_X1 \buffer_reg[14][1][0][2]  (.D(\input_filter[1][0] [2]), .CK(n_56_11), 
      .Q(\buffer[14][1][0] [2]), .QN());
   DFF_X1 \buffer_reg[14][1][0][1]  (.D(\input_filter[1][0] [1]), .CK(n_56_11), 
      .Q(\buffer[14][1][0] [1]), .QN());
   DFF_X1 \buffer_reg[14][1][0][0]  (.D(\input_filter[1][0] [0]), .CK(n_56_11), 
      .Q(\buffer[14][1][0] [0]), .QN());
   DFF_X1 \buffer_reg[13][1][0][15]  (.D(\input_filter[1][0] [15]), .CK(n_56_10), 
      .Q(\buffer[13][1][0] [15]), .QN());
   DFF_X1 \buffer_reg[13][1][0][14]  (.D(\input_filter[1][0] [14]), .CK(n_56_10), 
      .Q(\buffer[13][1][0] [14]), .QN());
   DFF_X1 \buffer_reg[13][1][0][13]  (.D(\input_filter[1][0] [13]), .CK(n_56_10), 
      .Q(\buffer[13][1][0] [13]), .QN());
   DFF_X1 \buffer_reg[13][1][0][12]  (.D(\input_filter[1][0] [12]), .CK(n_56_10), 
      .Q(\buffer[13][1][0] [12]), .QN());
   DFF_X1 \buffer_reg[13][1][0][11]  (.D(\input_filter[1][0] [11]), .CK(n_56_10), 
      .Q(\buffer[13][1][0] [11]), .QN());
   DFF_X1 \buffer_reg[13][1][0][10]  (.D(\input_filter[1][0] [10]), .CK(n_56_10), 
      .Q(\buffer[13][1][0] [10]), .QN());
   DFF_X1 \buffer_reg[13][1][0][9]  (.D(\input_filter[1][0] [9]), .CK(n_56_10), 
      .Q(\buffer[13][1][0] [9]), .QN());
   DFF_X1 \buffer_reg[13][1][0][8]  (.D(\input_filter[1][0] [8]), .CK(n_56_10), 
      .Q(\buffer[13][1][0] [8]), .QN());
   DFF_X1 \buffer_reg[13][1][0][7]  (.D(\input_filter[1][0] [7]), .CK(n_56_10), 
      .Q(\buffer[13][1][0] [7]), .QN());
   DFF_X1 \buffer_reg[13][1][0][6]  (.D(\input_filter[1][0] [6]), .CK(n_56_10), 
      .Q(\buffer[13][1][0] [6]), .QN());
   DFF_X1 \buffer_reg[13][1][0][5]  (.D(\input_filter[1][0] [5]), .CK(n_56_10), 
      .Q(\buffer[13][1][0] [5]), .QN());
   DFF_X1 \buffer_reg[13][1][0][4]  (.D(\input_filter[1][0] [4]), .CK(n_56_10), 
      .Q(\buffer[13][1][0] [4]), .QN());
   DFF_X1 \buffer_reg[13][1][0][3]  (.D(\input_filter[1][0] [3]), .CK(n_56_10), 
      .Q(\buffer[13][1][0] [3]), .QN());
   DFF_X1 \buffer_reg[13][1][0][2]  (.D(\input_filter[1][0] [2]), .CK(n_56_10), 
      .Q(\buffer[13][1][0] [2]), .QN());
   DFF_X1 \buffer_reg[13][1][0][1]  (.D(\input_filter[1][0] [1]), .CK(n_56_10), 
      .Q(\buffer[13][1][0] [1]), .QN());
   DFF_X1 \buffer_reg[13][1][0][0]  (.D(\input_filter[1][0] [0]), .CK(n_56_10), 
      .Q(\buffer[13][1][0] [0]), .QN());
   CLKGATETST_X1 \clk_gate_buffer_reg[3][0][0]_reg  (.CK(read), .E(n_3), 
      .SE(1'b0), .GCK(n_56_0));
   CLKGATETST_X1 \clk_gate_buffer_reg[4][0][0]_reg  (.CK(read), .E(n_4), 
      .SE(1'b0), .GCK(n_56_1));
   CLKGATETST_X1 \clk_gate_buffer_reg[5][0][0]_reg  (.CK(read), .E(n_5), 
      .SE(1'b0), .GCK(n_56_2));
   CLKGATETST_X1 \clk_gate_buffer_reg[6][0][0]_reg  (.CK(read), .E(n_6), 
      .SE(1'b0), .GCK(n_56_3));
   CLKGATETST_X1 \clk_gate_buffer_reg[7][0][0]_reg  (.CK(read), .E(n_7), 
      .SE(1'b0), .GCK(n_56_4));
   CLKGATETST_X1 \clk_gate_buffer_reg[8][0][0]_reg  (.CK(read), .E(n_8), 
      .SE(1'b0), .GCK(n_56_5));
   CLKGATETST_X1 \clk_gate_buffer_reg[9][0][0]_reg  (.CK(read), .E(n_9), 
      .SE(1'b0), .GCK(n_56_6));
   CLKGATETST_X1 \clk_gate_buffer_reg[10][0][0]_reg  (.CK(read), .E(n_10), 
      .SE(1'b0), .GCK(n_56_7));
   CLKGATETST_X1 \clk_gate_buffer_reg[11][0][0]_reg  (.CK(read), .E(n_11), 
      .SE(1'b0), .GCK(n_56_8));
   CLKGATETST_X1 \clk_gate_buffer_reg[12][0][0]_reg  (.CK(read), .E(n_12), 
      .SE(1'b0), .GCK(n_56_9));
   CLKGATETST_X1 \clk_gate_buffer_reg[13][0][0]_reg  (.CK(read), .E(n_13), 
      .SE(1'b0), .GCK(n_56_10));
   CLKGATETST_X1 \clk_gate_buffer_reg[14][0][0]_reg  (.CK(read), .E(n_14), 
      .SE(1'b0), .GCK(n_56_11));
   CLKGATETST_X1 \clk_gate_buffer_reg[0][0][1]_reg  (.CK(read), .E(n_0), 
      .SE(1'b0), .GCK(n_56_12));
   CLKGATETST_X1 \clk_gate_buffer_reg[1][0][1]_reg  (.CK(read), .E(n_1), 
      .SE(1'b0), .GCK(n_56_13));
   CLKGATETST_X1 \clk_gate_buffer_reg[2][0][1]_reg  (.CK(read), .E(n_2), 
      .SE(1'b0), .GCK(n_56_14));
   CLKGATETST_X1 \clk_gate_buffer_reg[15][0][1]_reg  (.CK(read), .E(n_15), 
      .SE(1'b0), .GCK(n_56_15));
   DFF_X1 \buffer_reg[0][1][2][15]  (.D(\input_filter[1][2] [15]), .CK(n_57_4), 
      .Q(\buffer[0][1][2] [15]), .QN());
   DFF_X1 \buffer_reg[0][1][2][14]  (.D(\input_filter[1][2] [14]), .CK(n_57_4), 
      .Q(\buffer[0][1][2] [14]), .QN());
   DFF_X1 \buffer_reg[0][1][2][13]  (.D(\input_filter[1][2] [13]), .CK(n_57_4), 
      .Q(\buffer[0][1][2] [13]), .QN());
   DFF_X1 \buffer_reg[0][1][2][12]  (.D(\input_filter[1][2] [12]), .CK(n_57_4), 
      .Q(\buffer[0][1][2] [12]), .QN());
   DFF_X1 \buffer_reg[0][1][2][11]  (.D(\input_filter[1][2] [11]), .CK(n_57_4), 
      .Q(\buffer[0][1][2] [11]), .QN());
   DFF_X1 \buffer_reg[0][1][2][10]  (.D(\input_filter[1][2] [10]), .CK(n_57_4), 
      .Q(\buffer[0][1][2] [10]), .QN());
   DFF_X1 \buffer_reg[0][1][2][9]  (.D(\input_filter[1][2] [9]), .CK(n_57_4), 
      .Q(\buffer[0][1][2] [9]), .QN());
   DFF_X1 \buffer_reg[0][1][2][8]  (.D(\input_filter[1][2] [8]), .CK(n_57_4), 
      .Q(\buffer[0][1][2] [8]), .QN());
   DFF_X1 \buffer_reg[0][1][2][7]  (.D(\input_filter[1][2] [7]), .CK(n_57_4), 
      .Q(\buffer[0][1][2] [7]), .QN());
   DFF_X1 \buffer_reg[0][1][2][6]  (.D(\input_filter[1][2] [6]), .CK(n_57_4), 
      .Q(\buffer[0][1][2] [6]), .QN());
   DFF_X1 \buffer_reg[0][1][2][5]  (.D(\input_filter[1][2] [5]), .CK(n_57_4), 
      .Q(\buffer[0][1][2] [5]), .QN());
   DFF_X1 \buffer_reg[0][1][2][4]  (.D(\input_filter[1][2] [4]), .CK(n_57_4), 
      .Q(\buffer[0][1][2] [4]), .QN());
   DFF_X1 \buffer_reg[0][1][2][3]  (.D(\input_filter[1][2] [3]), .CK(n_57_4), 
      .Q(\buffer[0][1][2] [3]), .QN());
   DFF_X1 \buffer_reg[0][1][2][2]  (.D(\input_filter[1][2] [2]), .CK(n_57_4), 
      .Q(\buffer[0][1][2] [2]), .QN());
   DFF_X1 \buffer_reg[0][1][2][1]  (.D(\input_filter[1][2] [1]), .CK(n_57_4), 
      .Q(\buffer[0][1][2] [1]), .QN());
   DFF_X1 \buffer_reg[0][1][2][0]  (.D(\input_filter[1][2] [0]), .CK(n_57_4), 
      .Q(\buffer[0][1][2] [0]), .QN());
   DFF_X1 \buffer_reg[9][1][2][15]  (.D(\input_filter[1][2] [15]), .CK(n_57_5), 
      .Q(\buffer[9][1][2] [15]), .QN());
   DFF_X1 \buffer_reg[9][1][2][14]  (.D(\input_filter[1][2] [14]), .CK(n_57_5), 
      .Q(\buffer[9][1][2] [14]), .QN());
   DFF_X1 \buffer_reg[9][1][2][13]  (.D(\input_filter[1][2] [13]), .CK(n_57_5), 
      .Q(\buffer[9][1][2] [13]), .QN());
   DFF_X1 \buffer_reg[9][1][2][12]  (.D(\input_filter[1][2] [12]), .CK(n_57_5), 
      .Q(\buffer[9][1][2] [12]), .QN());
   DFF_X1 \buffer_reg[9][1][2][11]  (.D(\input_filter[1][2] [11]), .CK(n_57_5), 
      .Q(\buffer[9][1][2] [11]), .QN());
   DFF_X1 \buffer_reg[9][1][2][10]  (.D(\input_filter[1][2] [10]), .CK(n_57_5), 
      .Q(\buffer[9][1][2] [10]), .QN());
   DFF_X1 \buffer_reg[9][1][2][9]  (.D(\input_filter[1][2] [9]), .CK(n_57_5), 
      .Q(\buffer[9][1][2] [9]), .QN());
   DFF_X1 \buffer_reg[9][1][2][8]  (.D(\input_filter[1][2] [8]), .CK(n_57_5), 
      .Q(\buffer[9][1][2] [8]), .QN());
   DFF_X1 \buffer_reg[9][1][2][7]  (.D(\input_filter[1][2] [7]), .CK(n_57_5), 
      .Q(\buffer[9][1][2] [7]), .QN());
   DFF_X1 \buffer_reg[9][1][2][6]  (.D(\input_filter[1][2] [6]), .CK(n_57_5), 
      .Q(\buffer[9][1][2] [6]), .QN());
   DFF_X1 \buffer_reg[9][1][2][5]  (.D(\input_filter[1][2] [5]), .CK(n_57_5), 
      .Q(\buffer[9][1][2] [5]), .QN());
   DFF_X1 \buffer_reg[9][1][2][4]  (.D(\input_filter[1][2] [4]), .CK(n_57_5), 
      .Q(\buffer[9][1][2] [4]), .QN());
   DFF_X1 \buffer_reg[9][1][2][3]  (.D(\input_filter[1][2] [3]), .CK(n_57_5), 
      .Q(\buffer[9][1][2] [3]), .QN());
   DFF_X1 \buffer_reg[9][1][2][2]  (.D(\input_filter[1][2] [2]), .CK(n_57_5), 
      .Q(\buffer[9][1][2] [2]), .QN());
   DFF_X1 \buffer_reg[9][1][2][1]  (.D(\input_filter[1][2] [1]), .CK(n_57_5), 
      .Q(\buffer[9][1][2] [1]), .QN());
   DFF_X1 \buffer_reg[9][1][2][0]  (.D(\input_filter[1][2] [0]), .CK(n_57_5), 
      .Q(\buffer[9][1][2] [0]), .QN());
   DFF_X1 \buffer_reg[10][1][2][15]  (.D(\input_filter[1][2] [15]), .CK(n_57_6), 
      .Q(\buffer[10][1][2] [15]), .QN());
   DFF_X1 \buffer_reg[10][1][2][14]  (.D(\input_filter[1][2] [14]), .CK(n_57_6), 
      .Q(\buffer[10][1][2] [14]), .QN());
   DFF_X1 \buffer_reg[10][1][2][13]  (.D(\input_filter[1][2] [13]), .CK(n_57_6), 
      .Q(\buffer[10][1][2] [13]), .QN());
   DFF_X1 \buffer_reg[10][1][2][12]  (.D(\input_filter[1][2] [12]), .CK(n_57_6), 
      .Q(\buffer[10][1][2] [12]), .QN());
   DFF_X1 \buffer_reg[10][1][2][11]  (.D(\input_filter[1][2] [11]), .CK(n_57_6), 
      .Q(\buffer[10][1][2] [11]), .QN());
   DFF_X1 \buffer_reg[10][1][2][10]  (.D(\input_filter[1][2] [10]), .CK(n_57_6), 
      .Q(\buffer[10][1][2] [10]), .QN());
   DFF_X1 \buffer_reg[10][1][2][9]  (.D(\input_filter[1][2] [9]), .CK(n_57_6), 
      .Q(\buffer[10][1][2] [9]), .QN());
   DFF_X1 \buffer_reg[10][1][2][8]  (.D(\input_filter[1][2] [8]), .CK(n_57_6), 
      .Q(\buffer[10][1][2] [8]), .QN());
   DFF_X1 \buffer_reg[10][1][2][7]  (.D(\input_filter[1][2] [7]), .CK(n_57_6), 
      .Q(\buffer[10][1][2] [7]), .QN());
   DFF_X1 \buffer_reg[10][1][2][6]  (.D(\input_filter[1][2] [6]), .CK(n_57_6), 
      .Q(\buffer[10][1][2] [6]), .QN());
   DFF_X1 \buffer_reg[10][1][2][5]  (.D(\input_filter[1][2] [5]), .CK(n_57_6), 
      .Q(\buffer[10][1][2] [5]), .QN());
   DFF_X1 \buffer_reg[10][1][2][4]  (.D(\input_filter[1][2] [4]), .CK(n_57_6), 
      .Q(\buffer[10][1][2] [4]), .QN());
   DFF_X1 \buffer_reg[10][1][2][3]  (.D(\input_filter[1][2] [3]), .CK(n_57_6), 
      .Q(\buffer[10][1][2] [3]), .QN());
   DFF_X1 \buffer_reg[10][1][2][2]  (.D(\input_filter[1][2] [2]), .CK(n_57_6), 
      .Q(\buffer[10][1][2] [2]), .QN());
   DFF_X1 \buffer_reg[10][1][2][1]  (.D(\input_filter[1][2] [1]), .CK(n_57_6), 
      .Q(\buffer[10][1][2] [1]), .QN());
   DFF_X1 \buffer_reg[10][1][2][0]  (.D(\input_filter[1][2] [0]), .CK(n_57_6), 
      .Q(\buffer[10][1][2] [0]), .QN());
   DFF_X1 \buffer_reg[11][1][2][15]  (.D(\input_filter[1][2] [15]), .CK(n_57_7), 
      .Q(\buffer[11][1][2] [15]), .QN());
   DFF_X1 \buffer_reg[11][1][2][14]  (.D(\input_filter[1][2] [14]), .CK(n_57_7), 
      .Q(\buffer[11][1][2] [14]), .QN());
   DFF_X1 \buffer_reg[11][1][2][13]  (.D(\input_filter[1][2] [13]), .CK(n_57_7), 
      .Q(\buffer[11][1][2] [13]), .QN());
   DFF_X1 \buffer_reg[11][1][2][12]  (.D(\input_filter[1][2] [12]), .CK(n_57_7), 
      .Q(\buffer[11][1][2] [12]), .QN());
   DFF_X1 \buffer_reg[11][1][2][11]  (.D(\input_filter[1][2] [11]), .CK(n_57_7), 
      .Q(\buffer[11][1][2] [11]), .QN());
   DFF_X1 \buffer_reg[11][1][2][10]  (.D(\input_filter[1][2] [10]), .CK(n_57_7), 
      .Q(\buffer[11][1][2] [10]), .QN());
   DFF_X1 \buffer_reg[11][1][2][9]  (.D(\input_filter[1][2] [9]), .CK(n_57_7), 
      .Q(\buffer[11][1][2] [9]), .QN());
   DFF_X1 \buffer_reg[11][1][2][8]  (.D(\input_filter[1][2] [8]), .CK(n_57_7), 
      .Q(\buffer[11][1][2] [8]), .QN());
   DFF_X1 \buffer_reg[11][1][2][7]  (.D(\input_filter[1][2] [7]), .CK(n_57_7), 
      .Q(\buffer[11][1][2] [7]), .QN());
   DFF_X1 \buffer_reg[11][1][2][6]  (.D(\input_filter[1][2] [6]), .CK(n_57_7), 
      .Q(\buffer[11][1][2] [6]), .QN());
   DFF_X1 \buffer_reg[11][1][2][5]  (.D(\input_filter[1][2] [5]), .CK(n_57_7), 
      .Q(\buffer[11][1][2] [5]), .QN());
   DFF_X1 \buffer_reg[11][1][2][4]  (.D(\input_filter[1][2] [4]), .CK(n_57_7), 
      .Q(\buffer[11][1][2] [4]), .QN());
   DFF_X1 \buffer_reg[11][1][2][3]  (.D(\input_filter[1][2] [3]), .CK(n_57_7), 
      .Q(\buffer[11][1][2] [3]), .QN());
   DFF_X1 \buffer_reg[11][1][2][2]  (.D(\input_filter[1][2] [2]), .CK(n_57_7), 
      .Q(\buffer[11][1][2] [2]), .QN());
   DFF_X1 \buffer_reg[11][1][2][1]  (.D(\input_filter[1][2] [1]), .CK(n_57_7), 
      .Q(\buffer[11][1][2] [1]), .QN());
   DFF_X1 \buffer_reg[11][1][2][0]  (.D(\input_filter[1][2] [0]), .CK(n_57_7), 
      .Q(\buffer[11][1][2] [0]), .QN());
   DFF_X1 \buffer_reg[12][1][2][15]  (.D(\input_filter[1][2] [15]), .CK(n_57_12), 
      .Q(\buffer[12][1][2] [15]), .QN());
   DFF_X1 \buffer_reg[12][1][2][14]  (.D(\input_filter[1][2] [14]), .CK(n_57_12), 
      .Q(\buffer[12][1][2] [14]), .QN());
   DFF_X1 \buffer_reg[12][1][2][13]  (.D(\input_filter[1][2] [13]), .CK(n_57_12), 
      .Q(\buffer[12][1][2] [13]), .QN());
   DFF_X1 \buffer_reg[12][1][2][12]  (.D(\input_filter[1][2] [12]), .CK(n_57_12), 
      .Q(\buffer[12][1][2] [12]), .QN());
   DFF_X1 \buffer_reg[12][1][2][11]  (.D(\input_filter[1][2] [11]), .CK(n_57_12), 
      .Q(\buffer[12][1][2] [11]), .QN());
   DFF_X1 \buffer_reg[12][1][2][10]  (.D(\input_filter[1][2] [10]), .CK(n_57_12), 
      .Q(\buffer[12][1][2] [10]), .QN());
   DFF_X1 \buffer_reg[12][1][2][9]  (.D(\input_filter[1][2] [9]), .CK(n_57_12), 
      .Q(\buffer[12][1][2] [9]), .QN());
   DFF_X1 \buffer_reg[12][1][2][8]  (.D(\input_filter[1][2] [8]), .CK(n_57_12), 
      .Q(\buffer[12][1][2] [8]), .QN());
   DFF_X1 \buffer_reg[12][1][2][7]  (.D(\input_filter[1][2] [7]), .CK(n_57_12), 
      .Q(\buffer[12][1][2] [7]), .QN());
   DFF_X1 \buffer_reg[12][1][2][6]  (.D(\input_filter[1][2] [6]), .CK(n_57_12), 
      .Q(\buffer[12][1][2] [6]), .QN());
   DFF_X1 \buffer_reg[12][1][2][5]  (.D(\input_filter[1][2] [5]), .CK(n_57_12), 
      .Q(\buffer[12][1][2] [5]), .QN());
   DFF_X1 \buffer_reg[12][1][2][4]  (.D(\input_filter[1][2] [4]), .CK(n_57_12), 
      .Q(\buffer[12][1][2] [4]), .QN());
   DFF_X1 \buffer_reg[12][1][2][3]  (.D(\input_filter[1][2] [3]), .CK(n_57_12), 
      .Q(\buffer[12][1][2] [3]), .QN());
   DFF_X1 \buffer_reg[12][1][2][2]  (.D(\input_filter[1][2] [2]), .CK(n_57_12), 
      .Q(\buffer[12][1][2] [2]), .QN());
   DFF_X1 \buffer_reg[12][1][2][1]  (.D(\input_filter[1][2] [1]), .CK(n_57_12), 
      .Q(\buffer[12][1][2] [1]), .QN());
   DFF_X1 \buffer_reg[12][1][2][0]  (.D(\input_filter[1][2] [0]), .CK(n_57_12), 
      .Q(\buffer[12][1][2] [0]), .QN());
   DFF_X1 \buffer_reg[13][1][2][15]  (.D(\input_filter[1][2] [15]), .CK(n_57_13), 
      .Q(\buffer[13][1][2] [15]), .QN());
   DFF_X1 \buffer_reg[13][1][2][14]  (.D(\input_filter[1][2] [14]), .CK(n_57_13), 
      .Q(\buffer[13][1][2] [14]), .QN());
   DFF_X1 \buffer_reg[13][1][2][13]  (.D(\input_filter[1][2] [13]), .CK(n_57_13), 
      .Q(\buffer[13][1][2] [13]), .QN());
   DFF_X1 \buffer_reg[13][1][2][12]  (.D(\input_filter[1][2] [12]), .CK(n_57_13), 
      .Q(\buffer[13][1][2] [12]), .QN());
   DFF_X1 \buffer_reg[13][1][2][11]  (.D(\input_filter[1][2] [11]), .CK(n_57_13), 
      .Q(\buffer[13][1][2] [11]), .QN());
   DFF_X1 \buffer_reg[13][1][2][10]  (.D(\input_filter[1][2] [10]), .CK(n_57_13), 
      .Q(\buffer[13][1][2] [10]), .QN());
   DFF_X1 \buffer_reg[13][1][2][9]  (.D(\input_filter[1][2] [9]), .CK(n_57_13), 
      .Q(\buffer[13][1][2] [9]), .QN());
   DFF_X1 \buffer_reg[13][1][2][8]  (.D(\input_filter[1][2] [8]), .CK(n_57_13), 
      .Q(\buffer[13][1][2] [8]), .QN());
   DFF_X1 \buffer_reg[13][1][2][7]  (.D(\input_filter[1][2] [7]), .CK(n_57_13), 
      .Q(\buffer[13][1][2] [7]), .QN());
   DFF_X1 \buffer_reg[13][1][2][6]  (.D(\input_filter[1][2] [6]), .CK(n_57_13), 
      .Q(\buffer[13][1][2] [6]), .QN());
   DFF_X1 \buffer_reg[13][1][2][5]  (.D(\input_filter[1][2] [5]), .CK(n_57_13), 
      .Q(\buffer[13][1][2] [5]), .QN());
   DFF_X1 \buffer_reg[13][1][2][4]  (.D(\input_filter[1][2] [4]), .CK(n_57_13), 
      .Q(\buffer[13][1][2] [4]), .QN());
   DFF_X1 \buffer_reg[13][1][2][3]  (.D(\input_filter[1][2] [3]), .CK(n_57_13), 
      .Q(\buffer[13][1][2] [3]), .QN());
   DFF_X1 \buffer_reg[13][1][2][2]  (.D(\input_filter[1][2] [2]), .CK(n_57_13), 
      .Q(\buffer[13][1][2] [2]), .QN());
   DFF_X1 \buffer_reg[13][1][2][1]  (.D(\input_filter[1][2] [1]), .CK(n_57_13), 
      .Q(\buffer[13][1][2] [1]), .QN());
   DFF_X1 \buffer_reg[13][1][2][0]  (.D(\input_filter[1][2] [0]), .CK(n_57_13), 
      .Q(\buffer[13][1][2] [0]), .QN());
   DFF_X1 \buffer_reg[14][1][2][15]  (.D(\input_filter[1][2] [15]), .CK(n_57_14), 
      .Q(\buffer[14][1][2] [15]), .QN());
   DFF_X1 \buffer_reg[14][1][2][14]  (.D(\input_filter[1][2] [14]), .CK(n_57_14), 
      .Q(\buffer[14][1][2] [14]), .QN());
   DFF_X1 \buffer_reg[14][1][2][13]  (.D(\input_filter[1][2] [13]), .CK(n_57_14), 
      .Q(\buffer[14][1][2] [13]), .QN());
   DFF_X1 \buffer_reg[14][1][2][12]  (.D(\input_filter[1][2] [12]), .CK(n_57_14), 
      .Q(\buffer[14][1][2] [12]), .QN());
   DFF_X1 \buffer_reg[14][1][2][11]  (.D(\input_filter[1][2] [11]), .CK(n_57_14), 
      .Q(\buffer[14][1][2] [11]), .QN());
   DFF_X1 \buffer_reg[14][1][2][10]  (.D(\input_filter[1][2] [10]), .CK(n_57_14), 
      .Q(\buffer[14][1][2] [10]), .QN());
   DFF_X1 \buffer_reg[14][1][2][9]  (.D(\input_filter[1][2] [9]), .CK(n_57_14), 
      .Q(\buffer[14][1][2] [9]), .QN());
   DFF_X1 \buffer_reg[14][1][2][8]  (.D(\input_filter[1][2] [8]), .CK(n_57_14), 
      .Q(\buffer[14][1][2] [8]), .QN());
   DFF_X1 \buffer_reg[14][1][2][7]  (.D(\input_filter[1][2] [7]), .CK(n_57_14), 
      .Q(\buffer[14][1][2] [7]), .QN());
   DFF_X1 \buffer_reg[14][1][2][6]  (.D(\input_filter[1][2] [6]), .CK(n_57_14), 
      .Q(\buffer[14][1][2] [6]), .QN());
   DFF_X1 \buffer_reg[14][1][2][5]  (.D(\input_filter[1][2] [5]), .CK(n_57_14), 
      .Q(\buffer[14][1][2] [5]), .QN());
   DFF_X1 \buffer_reg[14][1][2][4]  (.D(\input_filter[1][2] [4]), .CK(n_57_14), 
      .Q(\buffer[14][1][2] [4]), .QN());
   DFF_X1 \buffer_reg[14][1][2][3]  (.D(\input_filter[1][2] [3]), .CK(n_57_14), 
      .Q(\buffer[14][1][2] [3]), .QN());
   DFF_X1 \buffer_reg[14][1][2][2]  (.D(\input_filter[1][2] [2]), .CK(n_57_14), 
      .Q(\buffer[14][1][2] [2]), .QN());
   DFF_X1 \buffer_reg[14][1][2][1]  (.D(\input_filter[1][2] [1]), .CK(n_57_14), 
      .Q(\buffer[14][1][2] [1]), .QN());
   DFF_X1 \buffer_reg[14][1][2][0]  (.D(\input_filter[1][2] [0]), .CK(n_57_14), 
      .Q(\buffer[14][1][2] [0]), .QN());
   DFF_X1 \buffer_reg[15][1][2][15]  (.D(\input_filter[1][2] [15]), .CK(n_57_15), 
      .Q(\buffer[15][1][2] [15]), .QN());
   DFF_X1 \buffer_reg[15][1][2][14]  (.D(\input_filter[1][2] [14]), .CK(n_57_15), 
      .Q(\buffer[15][1][2] [14]), .QN());
   DFF_X1 \buffer_reg[15][1][2][13]  (.D(\input_filter[1][2] [13]), .CK(n_57_15), 
      .Q(\buffer[15][1][2] [13]), .QN());
   DFF_X1 \buffer_reg[15][1][2][12]  (.D(\input_filter[1][2] [12]), .CK(n_57_15), 
      .Q(\buffer[15][1][2] [12]), .QN());
   DFF_X1 \buffer_reg[15][1][2][11]  (.D(\input_filter[1][2] [11]), .CK(n_57_15), 
      .Q(\buffer[15][1][2] [11]), .QN());
   DFF_X1 \buffer_reg[15][1][2][10]  (.D(\input_filter[1][2] [10]), .CK(n_57_15), 
      .Q(\buffer[15][1][2] [10]), .QN());
   DFF_X1 \buffer_reg[15][1][2][9]  (.D(\input_filter[1][2] [9]), .CK(n_57_15), 
      .Q(\buffer[15][1][2] [9]), .QN());
   DFF_X1 \buffer_reg[15][1][2][8]  (.D(\input_filter[1][2] [8]), .CK(n_57_15), 
      .Q(\buffer[15][1][2] [8]), .QN());
   DFF_X1 \buffer_reg[15][1][2][7]  (.D(\input_filter[1][2] [7]), .CK(n_57_15), 
      .Q(\buffer[15][1][2] [7]), .QN());
   DFF_X1 \buffer_reg[15][1][2][6]  (.D(\input_filter[1][2] [6]), .CK(n_57_15), 
      .Q(\buffer[15][1][2] [6]), .QN());
   DFF_X1 \buffer_reg[15][1][2][5]  (.D(\input_filter[1][2] [5]), .CK(n_57_15), 
      .Q(\buffer[15][1][2] [5]), .QN());
   DFF_X1 \buffer_reg[15][1][2][4]  (.D(\input_filter[1][2] [4]), .CK(n_57_15), 
      .Q(\buffer[15][1][2] [4]), .QN());
   DFF_X1 \buffer_reg[15][1][2][3]  (.D(\input_filter[1][2] [3]), .CK(n_57_15), 
      .Q(\buffer[15][1][2] [3]), .QN());
   DFF_X1 \buffer_reg[15][1][2][2]  (.D(\input_filter[1][2] [2]), .CK(n_57_15), 
      .Q(\buffer[15][1][2] [2]), .QN());
   DFF_X1 \buffer_reg[15][1][2][1]  (.D(\input_filter[1][2] [1]), .CK(n_57_15), 
      .Q(\buffer[15][1][2] [1]), .QN());
   DFF_X1 \buffer_reg[15][1][2][0]  (.D(\input_filter[1][2] [0]), .CK(n_57_15), 
      .Q(\buffer[15][1][2] [0]), .QN());
   CLKGATETST_X1 \clk_gate_buffer_reg[4][0][4]_reg  (.CK(read), .E(n_4), 
      .SE(1'b0), .GCK(n_57_8));
   DFF_X1 \buffer_reg[4][0][4][15]  (.D(\input_filter[0][4] [15]), .CK(n_57_8), 
      .Q(\buffer[4][0][4] [15]), .QN());
   DFF_X1 \buffer_reg[4][0][4][14]  (.D(\input_filter[0][4] [14]), .CK(n_57_8), 
      .Q(\buffer[4][0][4] [14]), .QN());
   DFF_X1 \buffer_reg[4][0][4][13]  (.D(\input_filter[0][4] [13]), .CK(n_57_8), 
      .Q(\buffer[4][0][4] [13]), .QN());
   DFF_X1 \buffer_reg[4][0][4][12]  (.D(\input_filter[0][4] [12]), .CK(n_57_8), 
      .Q(\buffer[4][0][4] [12]), .QN());
   DFF_X1 \buffer_reg[4][0][4][11]  (.D(\input_filter[0][4] [11]), .CK(n_57_8), 
      .Q(\buffer[4][0][4] [11]), .QN());
   DFF_X1 \buffer_reg[4][0][4][10]  (.D(\input_filter[0][4] [10]), .CK(n_57_8), 
      .Q(\buffer[4][0][4] [10]), .QN());
   DFF_X1 \buffer_reg[4][0][4][9]  (.D(\input_filter[0][4] [9]), .CK(n_57_8), 
      .Q(\buffer[4][0][4] [9]), .QN());
   DFF_X1 \buffer_reg[4][0][4][8]  (.D(\input_filter[0][4] [8]), .CK(n_57_8), 
      .Q(\buffer[4][0][4] [8]), .QN());
   DFF_X1 \buffer_reg[4][0][4][7]  (.D(\input_filter[0][4] [7]), .CK(n_57_8), 
      .Q(\buffer[4][0][4] [7]), .QN());
   DFF_X1 \buffer_reg[4][0][4][6]  (.D(\input_filter[0][4] [6]), .CK(n_57_8), 
      .Q(\buffer[4][0][4] [6]), .QN());
   DFF_X1 \buffer_reg[4][0][4][5]  (.D(\input_filter[0][4] [5]), .CK(n_57_8), 
      .Q(\buffer[4][0][4] [5]), .QN());
   DFF_X1 \buffer_reg[4][0][4][4]  (.D(\input_filter[0][4] [4]), .CK(n_57_8), 
      .Q(\buffer[4][0][4] [4]), .QN());
   DFF_X1 \buffer_reg[4][0][4][3]  (.D(\input_filter[0][4] [3]), .CK(n_57_8), 
      .Q(\buffer[4][0][4] [3]), .QN());
   DFF_X1 \buffer_reg[4][0][4][2]  (.D(\input_filter[0][4] [2]), .CK(n_57_8), 
      .Q(\buffer[4][0][4] [2]), .QN());
   DFF_X1 \buffer_reg[4][0][4][1]  (.D(\input_filter[0][4] [1]), .CK(n_57_8), 
      .Q(\buffer[4][0][4] [1]), .QN());
   DFF_X1 \buffer_reg[4][0][4][0]  (.D(\input_filter[0][4] [0]), .CK(n_57_8), 
      .Q(\buffer[4][0][4] [0]), .QN());
   CLKGATETST_X1 \clk_gate_buffer_reg[3][0][4]_reg  (.CK(read), .E(n_3), 
      .SE(1'b0), .GCK(n_57_9));
   DFF_X1 \buffer_reg[3][0][4][15]  (.D(\input_filter[0][4] [15]), .CK(n_57_9), 
      .Q(\buffer[3][0][4] [15]), .QN());
   DFF_X1 \buffer_reg[3][0][4][14]  (.D(\input_filter[0][4] [14]), .CK(n_57_9), 
      .Q(\buffer[3][0][4] [14]), .QN());
   DFF_X1 \buffer_reg[3][0][4][13]  (.D(\input_filter[0][4] [13]), .CK(n_57_9), 
      .Q(\buffer[3][0][4] [13]), .QN());
   DFF_X1 \buffer_reg[3][0][4][12]  (.D(\input_filter[0][4] [12]), .CK(n_57_9), 
      .Q(\buffer[3][0][4] [12]), .QN());
   DFF_X1 \buffer_reg[3][0][4][11]  (.D(\input_filter[0][4] [11]), .CK(n_57_9), 
      .Q(\buffer[3][0][4] [11]), .QN());
   DFF_X1 \buffer_reg[3][0][4][10]  (.D(\input_filter[0][4] [10]), .CK(n_57_9), 
      .Q(\buffer[3][0][4] [10]), .QN());
   DFF_X1 \buffer_reg[3][0][4][9]  (.D(\input_filter[0][4] [9]), .CK(n_57_9), 
      .Q(\buffer[3][0][4] [9]), .QN());
   DFF_X1 \buffer_reg[3][0][4][8]  (.D(\input_filter[0][4] [8]), .CK(n_57_9), 
      .Q(\buffer[3][0][4] [8]), .QN());
   DFF_X1 \buffer_reg[3][0][4][7]  (.D(\input_filter[0][4] [7]), .CK(n_57_9), 
      .Q(\buffer[3][0][4] [7]), .QN());
   DFF_X1 \buffer_reg[3][0][4][6]  (.D(\input_filter[0][4] [6]), .CK(n_57_9), 
      .Q(\buffer[3][0][4] [6]), .QN());
   DFF_X1 \buffer_reg[3][0][4][5]  (.D(\input_filter[0][4] [5]), .CK(n_57_9), 
      .Q(\buffer[3][0][4] [5]), .QN());
   DFF_X1 \buffer_reg[3][0][4][4]  (.D(\input_filter[0][4] [4]), .CK(n_57_9), 
      .Q(\buffer[3][0][4] [4]), .QN());
   DFF_X1 \buffer_reg[3][0][4][3]  (.D(\input_filter[0][4] [3]), .CK(n_57_9), 
      .Q(\buffer[3][0][4] [3]), .QN());
   DFF_X1 \buffer_reg[3][0][4][2]  (.D(\input_filter[0][4] [2]), .CK(n_57_9), 
      .Q(\buffer[3][0][4] [2]), .QN());
   DFF_X1 \buffer_reg[3][0][4][1]  (.D(\input_filter[0][4] [1]), .CK(n_57_9), 
      .Q(\buffer[3][0][4] [1]), .QN());
   DFF_X1 \buffer_reg[3][0][4][0]  (.D(\input_filter[0][4] [0]), .CK(n_57_9), 
      .Q(\buffer[3][0][4] [0]), .QN());
   CLKGATETST_X1 \clk_gate_buffer_reg[2][0][4]_reg  (.CK(read), .E(n_2), 
      .SE(1'b0), .GCK(n_57_10));
   DFF_X1 \buffer_reg[2][0][4][15]  (.D(\input_filter[0][4] [15]), .CK(n_57_10), 
      .Q(\buffer[2][0][4] [15]), .QN());
   DFF_X1 \buffer_reg[2][0][4][14]  (.D(\input_filter[0][4] [14]), .CK(n_57_10), 
      .Q(\buffer[2][0][4] [14]), .QN());
   DFF_X1 \buffer_reg[2][0][4][13]  (.D(\input_filter[0][4] [13]), .CK(n_57_10), 
      .Q(\buffer[2][0][4] [13]), .QN());
   DFF_X1 \buffer_reg[2][0][4][12]  (.D(\input_filter[0][4] [12]), .CK(n_57_10), 
      .Q(\buffer[2][0][4] [12]), .QN());
   DFF_X1 \buffer_reg[2][0][4][11]  (.D(\input_filter[0][4] [11]), .CK(n_57_10), 
      .Q(\buffer[2][0][4] [11]), .QN());
   DFF_X1 \buffer_reg[2][0][4][10]  (.D(\input_filter[0][4] [10]), .CK(n_57_10), 
      .Q(\buffer[2][0][4] [10]), .QN());
   DFF_X1 \buffer_reg[2][0][4][9]  (.D(\input_filter[0][4] [9]), .CK(n_57_10), 
      .Q(\buffer[2][0][4] [9]), .QN());
   DFF_X1 \buffer_reg[2][0][4][8]  (.D(\input_filter[0][4] [8]), .CK(n_57_10), 
      .Q(\buffer[2][0][4] [8]), .QN());
   DFF_X1 \buffer_reg[2][0][4][7]  (.D(\input_filter[0][4] [7]), .CK(n_57_10), 
      .Q(\buffer[2][0][4] [7]), .QN());
   DFF_X1 \buffer_reg[2][0][4][6]  (.D(\input_filter[0][4] [6]), .CK(n_57_10), 
      .Q(\buffer[2][0][4] [6]), .QN());
   DFF_X1 \buffer_reg[2][0][4][5]  (.D(\input_filter[0][4] [5]), .CK(n_57_10), 
      .Q(\buffer[2][0][4] [5]), .QN());
   DFF_X1 \buffer_reg[2][0][4][4]  (.D(\input_filter[0][4] [4]), .CK(n_57_10), 
      .Q(\buffer[2][0][4] [4]), .QN());
   DFF_X1 \buffer_reg[2][0][4][3]  (.D(\input_filter[0][4] [3]), .CK(n_57_10), 
      .Q(\buffer[2][0][4] [3]), .QN());
   DFF_X1 \buffer_reg[2][0][4][2]  (.D(\input_filter[0][4] [2]), .CK(n_57_10), 
      .Q(\buffer[2][0][4] [2]), .QN());
   DFF_X1 \buffer_reg[2][0][4][1]  (.D(\input_filter[0][4] [1]), .CK(n_57_10), 
      .Q(\buffer[2][0][4] [1]), .QN());
   DFF_X1 \buffer_reg[2][0][4][0]  (.D(\input_filter[0][4] [0]), .CK(n_57_10), 
      .Q(\buffer[2][0][4] [0]), .QN());
   CLKGATETST_X1 \clk_gate_buffer_reg[1][0][4]_reg  (.CK(read), .E(n_1), 
      .SE(1'b0), .GCK(n_57_11));
   DFF_X1 \buffer_reg[1][0][4][15]  (.D(\input_filter[0][4] [15]), .CK(n_57_11), 
      .Q(\buffer[1][0][4] [15]), .QN());
   DFF_X1 \buffer_reg[1][0][4][14]  (.D(\input_filter[0][4] [14]), .CK(n_57_11), 
      .Q(\buffer[1][0][4] [14]), .QN());
   DFF_X1 \buffer_reg[1][0][4][13]  (.D(\input_filter[0][4] [13]), .CK(n_57_11), 
      .Q(\buffer[1][0][4] [13]), .QN());
   DFF_X1 \buffer_reg[1][0][4][12]  (.D(\input_filter[0][4] [12]), .CK(n_57_11), 
      .Q(\buffer[1][0][4] [12]), .QN());
   DFF_X1 \buffer_reg[1][0][4][11]  (.D(\input_filter[0][4] [11]), .CK(n_57_11), 
      .Q(\buffer[1][0][4] [11]), .QN());
   DFF_X1 \buffer_reg[1][0][4][10]  (.D(\input_filter[0][4] [10]), .CK(n_57_11), 
      .Q(\buffer[1][0][4] [10]), .QN());
   DFF_X1 \buffer_reg[1][0][4][9]  (.D(\input_filter[0][4] [9]), .CK(n_57_11), 
      .Q(\buffer[1][0][4] [9]), .QN());
   DFF_X1 \buffer_reg[1][0][4][8]  (.D(\input_filter[0][4] [8]), .CK(n_57_11), 
      .Q(\buffer[1][0][4] [8]), .QN());
   DFF_X1 \buffer_reg[1][0][4][7]  (.D(\input_filter[0][4] [7]), .CK(n_57_11), 
      .Q(\buffer[1][0][4] [7]), .QN());
   DFF_X1 \buffer_reg[1][0][4][6]  (.D(\input_filter[0][4] [6]), .CK(n_57_11), 
      .Q(\buffer[1][0][4] [6]), .QN());
   DFF_X1 \buffer_reg[1][0][4][5]  (.D(\input_filter[0][4] [5]), .CK(n_57_11), 
      .Q(\buffer[1][0][4] [5]), .QN());
   DFF_X1 \buffer_reg[1][0][4][4]  (.D(\input_filter[0][4] [4]), .CK(n_57_11), 
      .Q(\buffer[1][0][4] [4]), .QN());
   DFF_X1 \buffer_reg[1][0][4][3]  (.D(\input_filter[0][4] [3]), .CK(n_57_11), 
      .Q(\buffer[1][0][4] [3]), .QN());
   DFF_X1 \buffer_reg[1][0][4][2]  (.D(\input_filter[0][4] [2]), .CK(n_57_11), 
      .Q(\buffer[1][0][4] [2]), .QN());
   DFF_X1 \buffer_reg[1][0][4][1]  (.D(\input_filter[0][4] [1]), .CK(n_57_11), 
      .Q(\buffer[1][0][4] [1]), .QN());
   DFF_X1 \buffer_reg[1][0][4][0]  (.D(\input_filter[0][4] [0]), .CK(n_57_11), 
      .Q(\buffer[1][0][4] [0]), .QN());
   DFF_X1 \buffer_reg[0][0][4][15]  (.D(\input_filter[0][4] [15]), .CK(n_57_4), 
      .Q(\buffer[0][0][4] [15]), .QN());
   DFF_X1 \buffer_reg[0][0][4][14]  (.D(\input_filter[0][4] [14]), .CK(n_57_4), 
      .Q(\buffer[0][0][4] [14]), .QN());
   DFF_X1 \buffer_reg[0][0][4][13]  (.D(\input_filter[0][4] [13]), .CK(n_57_4), 
      .Q(\buffer[0][0][4] [13]), .QN());
   DFF_X1 \buffer_reg[0][0][4][12]  (.D(\input_filter[0][4] [12]), .CK(n_57_4), 
      .Q(\buffer[0][0][4] [12]), .QN());
   DFF_X1 \buffer_reg[0][0][4][11]  (.D(\input_filter[0][4] [11]), .CK(n_57_4), 
      .Q(\buffer[0][0][4] [11]), .QN());
   DFF_X1 \buffer_reg[0][0][4][10]  (.D(\input_filter[0][4] [10]), .CK(n_57_4), 
      .Q(\buffer[0][0][4] [10]), .QN());
   DFF_X1 \buffer_reg[0][0][4][9]  (.D(\input_filter[0][4] [9]), .CK(n_57_4), 
      .Q(\buffer[0][0][4] [9]), .QN());
   DFF_X1 \buffer_reg[0][0][4][8]  (.D(\input_filter[0][4] [8]), .CK(n_57_4), 
      .Q(\buffer[0][0][4] [8]), .QN());
   DFF_X1 \buffer_reg[0][0][4][7]  (.D(\input_filter[0][4] [7]), .CK(n_57_4), 
      .Q(\buffer[0][0][4] [7]), .QN());
   DFF_X1 \buffer_reg[0][0][4][6]  (.D(\input_filter[0][4] [6]), .CK(n_57_4), 
      .Q(\buffer[0][0][4] [6]), .QN());
   DFF_X1 \buffer_reg[0][0][4][5]  (.D(\input_filter[0][4] [5]), .CK(n_57_4), 
      .Q(\buffer[0][0][4] [5]), .QN());
   DFF_X1 \buffer_reg[0][0][4][4]  (.D(\input_filter[0][4] [4]), .CK(n_57_4), 
      .Q(\buffer[0][0][4] [4]), .QN());
   DFF_X1 \buffer_reg[0][0][4][3]  (.D(\input_filter[0][4] [3]), .CK(n_57_4), 
      .Q(\buffer[0][0][4] [3]), .QN());
   DFF_X1 \buffer_reg[0][0][4][2]  (.D(\input_filter[0][4] [2]), .CK(n_57_4), 
      .Q(\buffer[0][0][4] [2]), .QN());
   DFF_X1 \buffer_reg[0][0][4][1]  (.D(\input_filter[0][4] [1]), .CK(n_57_4), 
      .Q(\buffer[0][0][4] [1]), .QN());
   DFF_X1 \buffer_reg[0][0][4][0]  (.D(\input_filter[0][4] [0]), .CK(n_57_4), 
      .Q(\buffer[0][0][4] [0]), .QN());
   DFF_X1 \buffer_reg[15][0][4][15]  (.D(\input_filter[0][4] [15]), .CK(n_57_15), 
      .Q(\buffer[15][0][4] [15]), .QN());
   DFF_X1 \buffer_reg[15][0][4][14]  (.D(\input_filter[0][4] [14]), .CK(n_57_15), 
      .Q(\buffer[15][0][4] [14]), .QN());
   DFF_X1 \buffer_reg[15][0][4][13]  (.D(\input_filter[0][4] [13]), .CK(n_57_15), 
      .Q(\buffer[15][0][4] [13]), .QN());
   DFF_X1 \buffer_reg[15][0][4][12]  (.D(\input_filter[0][4] [12]), .CK(n_57_15), 
      .Q(\buffer[15][0][4] [12]), .QN());
   DFF_X1 \buffer_reg[15][0][4][11]  (.D(\input_filter[0][4] [11]), .CK(n_57_15), 
      .Q(\buffer[15][0][4] [11]), .QN());
   DFF_X1 \buffer_reg[15][0][4][10]  (.D(\input_filter[0][4] [10]), .CK(n_57_15), 
      .Q(\buffer[15][0][4] [10]), .QN());
   DFF_X1 \buffer_reg[15][0][4][9]  (.D(\input_filter[0][4] [9]), .CK(n_57_15), 
      .Q(\buffer[15][0][4] [9]), .QN());
   DFF_X1 \buffer_reg[15][0][4][8]  (.D(\input_filter[0][4] [8]), .CK(n_57_15), 
      .Q(\buffer[15][0][4] [8]), .QN());
   DFF_X1 \buffer_reg[15][0][4][7]  (.D(\input_filter[0][4] [7]), .CK(n_57_15), 
      .Q(\buffer[15][0][4] [7]), .QN());
   DFF_X1 \buffer_reg[15][0][4][6]  (.D(\input_filter[0][4] [6]), .CK(n_57_15), 
      .Q(\buffer[15][0][4] [6]), .QN());
   DFF_X1 \buffer_reg[15][0][4][5]  (.D(\input_filter[0][4] [5]), .CK(n_57_15), 
      .Q(\buffer[15][0][4] [5]), .QN());
   DFF_X1 \buffer_reg[15][0][4][4]  (.D(\input_filter[0][4] [4]), .CK(n_57_15), 
      .Q(\buffer[15][0][4] [4]), .QN());
   DFF_X1 \buffer_reg[15][0][4][3]  (.D(\input_filter[0][4] [3]), .CK(n_57_15), 
      .Q(\buffer[15][0][4] [3]), .QN());
   DFF_X1 \buffer_reg[15][0][4][2]  (.D(\input_filter[0][4] [2]), .CK(n_57_15), 
      .Q(\buffer[15][0][4] [2]), .QN());
   DFF_X1 \buffer_reg[15][0][4][1]  (.D(\input_filter[0][4] [1]), .CK(n_57_15), 
      .Q(\buffer[15][0][4] [1]), .QN());
   DFF_X1 \buffer_reg[15][0][4][0]  (.D(\input_filter[0][4] [0]), .CK(n_57_15), 
      .Q(\buffer[15][0][4] [0]), .QN());
   DFF_X1 \buffer_reg[14][0][4][15]  (.D(\input_filter[0][4] [15]), .CK(n_57_14), 
      .Q(\buffer[14][0][4] [15]), .QN());
   DFF_X1 \buffer_reg[14][0][4][14]  (.D(\input_filter[0][4] [14]), .CK(n_57_14), 
      .Q(\buffer[14][0][4] [14]), .QN());
   DFF_X1 \buffer_reg[14][0][4][13]  (.D(\input_filter[0][4] [13]), .CK(n_57_14), 
      .Q(\buffer[14][0][4] [13]), .QN());
   DFF_X1 \buffer_reg[14][0][4][12]  (.D(\input_filter[0][4] [12]), .CK(n_57_14), 
      .Q(\buffer[14][0][4] [12]), .QN());
   DFF_X1 \buffer_reg[14][0][4][11]  (.D(\input_filter[0][4] [11]), .CK(n_57_14), 
      .Q(\buffer[14][0][4] [11]), .QN());
   DFF_X1 \buffer_reg[14][0][4][10]  (.D(\input_filter[0][4] [10]), .CK(n_57_14), 
      .Q(\buffer[14][0][4] [10]), .QN());
   DFF_X1 \buffer_reg[14][0][4][9]  (.D(\input_filter[0][4] [9]), .CK(n_57_14), 
      .Q(\buffer[14][0][4] [9]), .QN());
   DFF_X1 \buffer_reg[14][0][4][8]  (.D(\input_filter[0][4] [8]), .CK(n_57_14), 
      .Q(\buffer[14][0][4] [8]), .QN());
   DFF_X1 \buffer_reg[14][0][4][7]  (.D(\input_filter[0][4] [7]), .CK(n_57_14), 
      .Q(\buffer[14][0][4] [7]), .QN());
   DFF_X1 \buffer_reg[14][0][4][6]  (.D(\input_filter[0][4] [6]), .CK(n_57_14), 
      .Q(\buffer[14][0][4] [6]), .QN());
   DFF_X1 \buffer_reg[14][0][4][5]  (.D(\input_filter[0][4] [5]), .CK(n_57_14), 
      .Q(\buffer[14][0][4] [5]), .QN());
   DFF_X1 \buffer_reg[14][0][4][4]  (.D(\input_filter[0][4] [4]), .CK(n_57_14), 
      .Q(\buffer[14][0][4] [4]), .QN());
   DFF_X1 \buffer_reg[14][0][4][3]  (.D(\input_filter[0][4] [3]), .CK(n_57_14), 
      .Q(\buffer[14][0][4] [3]), .QN());
   DFF_X1 \buffer_reg[14][0][4][2]  (.D(\input_filter[0][4] [2]), .CK(n_57_14), 
      .Q(\buffer[14][0][4] [2]), .QN());
   DFF_X1 \buffer_reg[14][0][4][1]  (.D(\input_filter[0][4] [1]), .CK(n_57_14), 
      .Q(\buffer[14][0][4] [1]), .QN());
   DFF_X1 \buffer_reg[14][0][4][0]  (.D(\input_filter[0][4] [0]), .CK(n_57_14), 
      .Q(\buffer[14][0][4] [0]), .QN());
   DFF_X1 \buffer_reg[13][0][4][15]  (.D(\input_filter[0][4] [15]), .CK(n_57_13), 
      .Q(\buffer[13][0][4] [15]), .QN());
   DFF_X1 \buffer_reg[13][0][4][14]  (.D(\input_filter[0][4] [14]), .CK(n_57_13), 
      .Q(\buffer[13][0][4] [14]), .QN());
   DFF_X1 \buffer_reg[13][0][4][13]  (.D(\input_filter[0][4] [13]), .CK(n_57_13), 
      .Q(\buffer[13][0][4] [13]), .QN());
   DFF_X1 \buffer_reg[13][0][4][12]  (.D(\input_filter[0][4] [12]), .CK(n_57_13), 
      .Q(\buffer[13][0][4] [12]), .QN());
   DFF_X1 \buffer_reg[13][0][4][11]  (.D(\input_filter[0][4] [11]), .CK(n_57_13), 
      .Q(\buffer[13][0][4] [11]), .QN());
   DFF_X1 \buffer_reg[13][0][4][10]  (.D(\input_filter[0][4] [10]), .CK(n_57_13), 
      .Q(\buffer[13][0][4] [10]), .QN());
   DFF_X1 \buffer_reg[13][0][4][9]  (.D(\input_filter[0][4] [9]), .CK(n_57_13), 
      .Q(\buffer[13][0][4] [9]), .QN());
   DFF_X1 \buffer_reg[13][0][4][8]  (.D(\input_filter[0][4] [8]), .CK(n_57_13), 
      .Q(\buffer[13][0][4] [8]), .QN());
   DFF_X1 \buffer_reg[13][0][4][7]  (.D(\input_filter[0][4] [7]), .CK(n_57_13), 
      .Q(\buffer[13][0][4] [7]), .QN());
   DFF_X1 \buffer_reg[13][0][4][6]  (.D(\input_filter[0][4] [6]), .CK(n_57_13), 
      .Q(\buffer[13][0][4] [6]), .QN());
   DFF_X1 \buffer_reg[13][0][4][5]  (.D(\input_filter[0][4] [5]), .CK(n_57_13), 
      .Q(\buffer[13][0][4] [5]), .QN());
   DFF_X1 \buffer_reg[13][0][4][4]  (.D(\input_filter[0][4] [4]), .CK(n_57_13), 
      .Q(\buffer[13][0][4] [4]), .QN());
   DFF_X1 \buffer_reg[13][0][4][3]  (.D(\input_filter[0][4] [3]), .CK(n_57_13), 
      .Q(\buffer[13][0][4] [3]), .QN());
   DFF_X1 \buffer_reg[13][0][4][2]  (.D(\input_filter[0][4] [2]), .CK(n_57_13), 
      .Q(\buffer[13][0][4] [2]), .QN());
   DFF_X1 \buffer_reg[13][0][4][1]  (.D(\input_filter[0][4] [1]), .CK(n_57_13), 
      .Q(\buffer[13][0][4] [1]), .QN());
   DFF_X1 \buffer_reg[13][0][4][0]  (.D(\input_filter[0][4] [0]), .CK(n_57_13), 
      .Q(\buffer[13][0][4] [0]), .QN());
   DFF_X1 \buffer_reg[12][0][4][15]  (.D(\input_filter[0][4] [15]), .CK(n_57_12), 
      .Q(\buffer[12][0][4] [15]), .QN());
   DFF_X1 \buffer_reg[12][0][4][14]  (.D(\input_filter[0][4] [14]), .CK(n_57_12), 
      .Q(\buffer[12][0][4] [14]), .QN());
   DFF_X1 \buffer_reg[12][0][4][13]  (.D(\input_filter[0][4] [13]), .CK(n_57_12), 
      .Q(\buffer[12][0][4] [13]), .QN());
   DFF_X1 \buffer_reg[12][0][4][12]  (.D(\input_filter[0][4] [12]), .CK(n_57_12), 
      .Q(\buffer[12][0][4] [12]), .QN());
   DFF_X1 \buffer_reg[12][0][4][11]  (.D(\input_filter[0][4] [11]), .CK(n_57_12), 
      .Q(\buffer[12][0][4] [11]), .QN());
   DFF_X1 \buffer_reg[12][0][4][10]  (.D(\input_filter[0][4] [10]), .CK(n_57_12), 
      .Q(\buffer[12][0][4] [10]), .QN());
   DFF_X1 \buffer_reg[12][0][4][9]  (.D(\input_filter[0][4] [9]), .CK(n_57_12), 
      .Q(\buffer[12][0][4] [9]), .QN());
   DFF_X1 \buffer_reg[12][0][4][8]  (.D(\input_filter[0][4] [8]), .CK(n_57_12), 
      .Q(\buffer[12][0][4] [8]), .QN());
   DFF_X1 \buffer_reg[12][0][4][7]  (.D(\input_filter[0][4] [7]), .CK(n_57_12), 
      .Q(\buffer[12][0][4] [7]), .QN());
   DFF_X1 \buffer_reg[12][0][4][6]  (.D(\input_filter[0][4] [6]), .CK(n_57_12), 
      .Q(\buffer[12][0][4] [6]), .QN());
   DFF_X1 \buffer_reg[12][0][4][5]  (.D(\input_filter[0][4] [5]), .CK(n_57_12), 
      .Q(\buffer[12][0][4] [5]), .QN());
   DFF_X1 \buffer_reg[12][0][4][4]  (.D(\input_filter[0][4] [4]), .CK(n_57_12), 
      .Q(\buffer[12][0][4] [4]), .QN());
   DFF_X1 \buffer_reg[12][0][4][3]  (.D(\input_filter[0][4] [3]), .CK(n_57_12), 
      .Q(\buffer[12][0][4] [3]), .QN());
   DFF_X1 \buffer_reg[12][0][4][2]  (.D(\input_filter[0][4] [2]), .CK(n_57_12), 
      .Q(\buffer[12][0][4] [2]), .QN());
   DFF_X1 \buffer_reg[12][0][4][1]  (.D(\input_filter[0][4] [1]), .CK(n_57_12), 
      .Q(\buffer[12][0][4] [1]), .QN());
   DFF_X1 \buffer_reg[12][0][4][0]  (.D(\input_filter[0][4] [0]), .CK(n_57_12), 
      .Q(\buffer[12][0][4] [0]), .QN());
   DFF_X1 \buffer_reg[11][0][4][15]  (.D(\input_filter[0][4] [15]), .CK(n_57_7), 
      .Q(\buffer[11][0][4] [15]), .QN());
   DFF_X1 \buffer_reg[11][0][4][14]  (.D(\input_filter[0][4] [14]), .CK(n_57_7), 
      .Q(\buffer[11][0][4] [14]), .QN());
   DFF_X1 \buffer_reg[11][0][4][13]  (.D(\input_filter[0][4] [13]), .CK(n_57_7), 
      .Q(\buffer[11][0][4] [13]), .QN());
   DFF_X1 \buffer_reg[11][0][4][12]  (.D(\input_filter[0][4] [12]), .CK(n_57_7), 
      .Q(\buffer[11][0][4] [12]), .QN());
   DFF_X1 \buffer_reg[11][0][4][11]  (.D(\input_filter[0][4] [11]), .CK(n_57_7), 
      .Q(\buffer[11][0][4] [11]), .QN());
   DFF_X1 \buffer_reg[11][0][4][10]  (.D(\input_filter[0][4] [10]), .CK(n_57_7), 
      .Q(\buffer[11][0][4] [10]), .QN());
   DFF_X1 \buffer_reg[11][0][4][9]  (.D(\input_filter[0][4] [9]), .CK(n_57_7), 
      .Q(\buffer[11][0][4] [9]), .QN());
   DFF_X1 \buffer_reg[11][0][4][8]  (.D(\input_filter[0][4] [8]), .CK(n_57_7), 
      .Q(\buffer[11][0][4] [8]), .QN());
   DFF_X1 \buffer_reg[11][0][4][7]  (.D(\input_filter[0][4] [7]), .CK(n_57_7), 
      .Q(\buffer[11][0][4] [7]), .QN());
   DFF_X1 \buffer_reg[11][0][4][6]  (.D(\input_filter[0][4] [6]), .CK(n_57_7), 
      .Q(\buffer[11][0][4] [6]), .QN());
   DFF_X1 \buffer_reg[11][0][4][5]  (.D(\input_filter[0][4] [5]), .CK(n_57_7), 
      .Q(\buffer[11][0][4] [5]), .QN());
   DFF_X1 \buffer_reg[11][0][4][4]  (.D(\input_filter[0][4] [4]), .CK(n_57_7), 
      .Q(\buffer[11][0][4] [4]), .QN());
   DFF_X1 \buffer_reg[11][0][4][3]  (.D(\input_filter[0][4] [3]), .CK(n_57_7), 
      .Q(\buffer[11][0][4] [3]), .QN());
   DFF_X1 \buffer_reg[11][0][4][2]  (.D(\input_filter[0][4] [2]), .CK(n_57_7), 
      .Q(\buffer[11][0][4] [2]), .QN());
   DFF_X1 \buffer_reg[11][0][4][1]  (.D(\input_filter[0][4] [1]), .CK(n_57_7), 
      .Q(\buffer[11][0][4] [1]), .QN());
   DFF_X1 \buffer_reg[11][0][4][0]  (.D(\input_filter[0][4] [0]), .CK(n_57_7), 
      .Q(\buffer[11][0][4] [0]), .QN());
   DFF_X1 \buffer_reg[10][0][4][15]  (.D(\input_filter[0][4] [15]), .CK(n_57_6), 
      .Q(\buffer[10][0][4] [15]), .QN());
   DFF_X1 \buffer_reg[10][0][4][14]  (.D(\input_filter[0][4] [14]), .CK(n_57_6), 
      .Q(\buffer[10][0][4] [14]), .QN());
   DFF_X1 \buffer_reg[10][0][4][13]  (.D(\input_filter[0][4] [13]), .CK(n_57_6), 
      .Q(\buffer[10][0][4] [13]), .QN());
   DFF_X1 \buffer_reg[10][0][4][12]  (.D(\input_filter[0][4] [12]), .CK(n_57_6), 
      .Q(\buffer[10][0][4] [12]), .QN());
   DFF_X1 \buffer_reg[10][0][4][11]  (.D(\input_filter[0][4] [11]), .CK(n_57_6), 
      .Q(\buffer[10][0][4] [11]), .QN());
   DFF_X1 \buffer_reg[10][0][4][10]  (.D(\input_filter[0][4] [10]), .CK(n_57_6), 
      .Q(\buffer[10][0][4] [10]), .QN());
   DFF_X1 \buffer_reg[10][0][4][9]  (.D(\input_filter[0][4] [9]), .CK(n_57_6), 
      .Q(\buffer[10][0][4] [9]), .QN());
   DFF_X1 \buffer_reg[10][0][4][8]  (.D(\input_filter[0][4] [8]), .CK(n_57_6), 
      .Q(\buffer[10][0][4] [8]), .QN());
   DFF_X1 \buffer_reg[10][0][4][7]  (.D(\input_filter[0][4] [7]), .CK(n_57_6), 
      .Q(\buffer[10][0][4] [7]), .QN());
   DFF_X1 \buffer_reg[10][0][4][6]  (.D(\input_filter[0][4] [6]), .CK(n_57_6), 
      .Q(\buffer[10][0][4] [6]), .QN());
   DFF_X1 \buffer_reg[10][0][4][5]  (.D(\input_filter[0][4] [5]), .CK(n_57_6), 
      .Q(\buffer[10][0][4] [5]), .QN());
   DFF_X1 \buffer_reg[10][0][4][4]  (.D(\input_filter[0][4] [4]), .CK(n_57_6), 
      .Q(\buffer[10][0][4] [4]), .QN());
   DFF_X1 \buffer_reg[10][0][4][3]  (.D(\input_filter[0][4] [3]), .CK(n_57_6), 
      .Q(\buffer[10][0][4] [3]), .QN());
   DFF_X1 \buffer_reg[10][0][4][2]  (.D(\input_filter[0][4] [2]), .CK(n_57_6), 
      .Q(\buffer[10][0][4] [2]), .QN());
   DFF_X1 \buffer_reg[10][0][4][1]  (.D(\input_filter[0][4] [1]), .CK(n_57_6), 
      .Q(\buffer[10][0][4] [1]), .QN());
   DFF_X1 \buffer_reg[10][0][4][0]  (.D(\input_filter[0][4] [0]), .CK(n_57_6), 
      .Q(\buffer[10][0][4] [0]), .QN());
   DFF_X1 \buffer_reg[9][0][4][15]  (.D(\input_filter[0][4] [15]), .CK(n_57_5), 
      .Q(\buffer[9][0][4] [15]), .QN());
   DFF_X1 \buffer_reg[9][0][4][14]  (.D(\input_filter[0][4] [14]), .CK(n_57_5), 
      .Q(\buffer[9][0][4] [14]), .QN());
   DFF_X1 \buffer_reg[9][0][4][13]  (.D(\input_filter[0][4] [13]), .CK(n_57_5), 
      .Q(\buffer[9][0][4] [13]), .QN());
   DFF_X1 \buffer_reg[9][0][4][12]  (.D(\input_filter[0][4] [12]), .CK(n_57_5), 
      .Q(\buffer[9][0][4] [12]), .QN());
   DFF_X1 \buffer_reg[9][0][4][11]  (.D(\input_filter[0][4] [11]), .CK(n_57_5), 
      .Q(\buffer[9][0][4] [11]), .QN());
   DFF_X1 \buffer_reg[9][0][4][10]  (.D(\input_filter[0][4] [10]), .CK(n_57_5), 
      .Q(\buffer[9][0][4] [10]), .QN());
   DFF_X1 \buffer_reg[9][0][4][9]  (.D(\input_filter[0][4] [9]), .CK(n_57_5), 
      .Q(\buffer[9][0][4] [9]), .QN());
   DFF_X1 \buffer_reg[9][0][4][8]  (.D(\input_filter[0][4] [8]), .CK(n_57_5), 
      .Q(\buffer[9][0][4] [8]), .QN());
   DFF_X1 \buffer_reg[9][0][4][7]  (.D(\input_filter[0][4] [7]), .CK(n_57_5), 
      .Q(\buffer[9][0][4] [7]), .QN());
   DFF_X1 \buffer_reg[9][0][4][6]  (.D(\input_filter[0][4] [6]), .CK(n_57_5), 
      .Q(\buffer[9][0][4] [6]), .QN());
   DFF_X1 \buffer_reg[9][0][4][5]  (.D(\input_filter[0][4] [5]), .CK(n_57_5), 
      .Q(\buffer[9][0][4] [5]), .QN());
   DFF_X1 \buffer_reg[9][0][4][4]  (.D(\input_filter[0][4] [4]), .CK(n_57_5), 
      .Q(\buffer[9][0][4] [4]), .QN());
   DFF_X1 \buffer_reg[9][0][4][3]  (.D(\input_filter[0][4] [3]), .CK(n_57_5), 
      .Q(\buffer[9][0][4] [3]), .QN());
   DFF_X1 \buffer_reg[9][0][4][2]  (.D(\input_filter[0][4] [2]), .CK(n_57_5), 
      .Q(\buffer[9][0][4] [2]), .QN());
   DFF_X1 \buffer_reg[9][0][4][1]  (.D(\input_filter[0][4] [1]), .CK(n_57_5), 
      .Q(\buffer[9][0][4] [1]), .QN());
   DFF_X1 \buffer_reg[9][0][4][0]  (.D(\input_filter[0][4] [0]), .CK(n_57_5), 
      .Q(\buffer[9][0][4] [0]), .QN());
   CLKGATETST_X1 \clk_gate_buffer_reg[8][0][4]_reg  (.CK(read), .E(n_8), 
      .SE(1'b0), .GCK(n_57_0));
   DFF_X1 \buffer_reg[8][0][4][15]  (.D(\input_filter[0][4] [15]), .CK(n_57_0), 
      .Q(\buffer[8][0][4] [15]), .QN());
   DFF_X1 \buffer_reg[8][0][4][14]  (.D(\input_filter[0][4] [14]), .CK(n_57_0), 
      .Q(\buffer[8][0][4] [14]), .QN());
   DFF_X1 \buffer_reg[8][0][4][13]  (.D(\input_filter[0][4] [13]), .CK(n_57_0), 
      .Q(\buffer[8][0][4] [13]), .QN());
   DFF_X1 \buffer_reg[8][0][4][12]  (.D(\input_filter[0][4] [12]), .CK(n_57_0), 
      .Q(\buffer[8][0][4] [12]), .QN());
   DFF_X1 \buffer_reg[8][0][4][11]  (.D(\input_filter[0][4] [11]), .CK(n_57_0), 
      .Q(\buffer[8][0][4] [11]), .QN());
   DFF_X1 \buffer_reg[8][0][4][10]  (.D(\input_filter[0][4] [10]), .CK(n_57_0), 
      .Q(\buffer[8][0][4] [10]), .QN());
   DFF_X1 \buffer_reg[8][0][4][9]  (.D(\input_filter[0][4] [9]), .CK(n_57_0), 
      .Q(\buffer[8][0][4] [9]), .QN());
   DFF_X1 \buffer_reg[8][0][4][8]  (.D(\input_filter[0][4] [8]), .CK(n_57_0), 
      .Q(\buffer[8][0][4] [8]), .QN());
   DFF_X1 \buffer_reg[8][0][4][7]  (.D(\input_filter[0][4] [7]), .CK(n_57_0), 
      .Q(\buffer[8][0][4] [7]), .QN());
   DFF_X1 \buffer_reg[8][0][4][6]  (.D(\input_filter[0][4] [6]), .CK(n_57_0), 
      .Q(\buffer[8][0][4] [6]), .QN());
   DFF_X1 \buffer_reg[8][0][4][5]  (.D(\input_filter[0][4] [5]), .CK(n_57_0), 
      .Q(\buffer[8][0][4] [5]), .QN());
   DFF_X1 \buffer_reg[8][0][4][4]  (.D(\input_filter[0][4] [4]), .CK(n_57_0), 
      .Q(\buffer[8][0][4] [4]), .QN());
   DFF_X1 \buffer_reg[8][0][4][3]  (.D(\input_filter[0][4] [3]), .CK(n_57_0), 
      .Q(\buffer[8][0][4] [3]), .QN());
   DFF_X1 \buffer_reg[8][0][4][2]  (.D(\input_filter[0][4] [2]), .CK(n_57_0), 
      .Q(\buffer[8][0][4] [2]), .QN());
   DFF_X1 \buffer_reg[8][0][4][1]  (.D(\input_filter[0][4] [1]), .CK(n_57_0), 
      .Q(\buffer[8][0][4] [1]), .QN());
   DFF_X1 \buffer_reg[8][0][4][0]  (.D(\input_filter[0][4] [0]), .CK(n_57_0), 
      .Q(\buffer[8][0][4] [0]), .QN());
   CLKGATETST_X1 \clk_gate_buffer_reg[7][0][4]_reg  (.CK(read), .E(n_7), 
      .SE(1'b0), .GCK(n_57_1));
   DFF_X1 \buffer_reg[7][0][4][15]  (.D(\input_filter[0][4] [15]), .CK(n_57_1), 
      .Q(\buffer[7][0][4] [15]), .QN());
   DFF_X1 \buffer_reg[7][0][4][14]  (.D(\input_filter[0][4] [14]), .CK(n_57_1), 
      .Q(\buffer[7][0][4] [14]), .QN());
   DFF_X1 \buffer_reg[7][0][4][13]  (.D(\input_filter[0][4] [13]), .CK(n_57_1), 
      .Q(\buffer[7][0][4] [13]), .QN());
   DFF_X1 \buffer_reg[7][0][4][12]  (.D(\input_filter[0][4] [12]), .CK(n_57_1), 
      .Q(\buffer[7][0][4] [12]), .QN());
   DFF_X1 \buffer_reg[7][0][4][11]  (.D(\input_filter[0][4] [11]), .CK(n_57_1), 
      .Q(\buffer[7][0][4] [11]), .QN());
   DFF_X1 \buffer_reg[7][0][4][10]  (.D(\input_filter[0][4] [10]), .CK(n_57_1), 
      .Q(\buffer[7][0][4] [10]), .QN());
   DFF_X1 \buffer_reg[7][0][4][9]  (.D(\input_filter[0][4] [9]), .CK(n_57_1), 
      .Q(\buffer[7][0][4] [9]), .QN());
   DFF_X1 \buffer_reg[7][0][4][8]  (.D(\input_filter[0][4] [8]), .CK(n_57_1), 
      .Q(\buffer[7][0][4] [8]), .QN());
   DFF_X1 \buffer_reg[7][0][4][7]  (.D(\input_filter[0][4] [7]), .CK(n_57_1), 
      .Q(\buffer[7][0][4] [7]), .QN());
   DFF_X1 \buffer_reg[7][0][4][6]  (.D(\input_filter[0][4] [6]), .CK(n_57_1), 
      .Q(\buffer[7][0][4] [6]), .QN());
   DFF_X1 \buffer_reg[7][0][4][5]  (.D(\input_filter[0][4] [5]), .CK(n_57_1), 
      .Q(\buffer[7][0][4] [5]), .QN());
   DFF_X1 \buffer_reg[7][0][4][4]  (.D(\input_filter[0][4] [4]), .CK(n_57_1), 
      .Q(\buffer[7][0][4] [4]), .QN());
   DFF_X1 \buffer_reg[7][0][4][3]  (.D(\input_filter[0][4] [3]), .CK(n_57_1), 
      .Q(\buffer[7][0][4] [3]), .QN());
   DFF_X1 \buffer_reg[7][0][4][2]  (.D(\input_filter[0][4] [2]), .CK(n_57_1), 
      .Q(\buffer[7][0][4] [2]), .QN());
   DFF_X1 \buffer_reg[7][0][4][1]  (.D(\input_filter[0][4] [1]), .CK(n_57_1), 
      .Q(\buffer[7][0][4] [1]), .QN());
   DFF_X1 \buffer_reg[7][0][4][0]  (.D(\input_filter[0][4] [0]), .CK(n_57_1), 
      .Q(\buffer[7][0][4] [0]), .QN());
   CLKGATETST_X1 \clk_gate_buffer_reg[6][0][4]_reg  (.CK(read), .E(n_6), 
      .SE(1'b0), .GCK(n_57_2));
   DFF_X1 \buffer_reg[6][0][4][15]  (.D(\input_filter[0][4] [15]), .CK(n_57_2), 
      .Q(\buffer[6][0][4] [15]), .QN());
   DFF_X1 \buffer_reg[6][0][4][14]  (.D(\input_filter[0][4] [14]), .CK(n_57_2), 
      .Q(\buffer[6][0][4] [14]), .QN());
   DFF_X1 \buffer_reg[6][0][4][13]  (.D(\input_filter[0][4] [13]), .CK(n_57_2), 
      .Q(\buffer[6][0][4] [13]), .QN());
   DFF_X1 \buffer_reg[6][0][4][12]  (.D(\input_filter[0][4] [12]), .CK(n_57_2), 
      .Q(\buffer[6][0][4] [12]), .QN());
   DFF_X1 \buffer_reg[6][0][4][11]  (.D(\input_filter[0][4] [11]), .CK(n_57_2), 
      .Q(\buffer[6][0][4] [11]), .QN());
   DFF_X1 \buffer_reg[6][0][4][10]  (.D(\input_filter[0][4] [10]), .CK(n_57_2), 
      .Q(\buffer[6][0][4] [10]), .QN());
   DFF_X1 \buffer_reg[6][0][4][9]  (.D(\input_filter[0][4] [9]), .CK(n_57_2), 
      .Q(\buffer[6][0][4] [9]), .QN());
   DFF_X1 \buffer_reg[6][0][4][8]  (.D(\input_filter[0][4] [8]), .CK(n_57_2), 
      .Q(\buffer[6][0][4] [8]), .QN());
   DFF_X1 \buffer_reg[6][0][4][7]  (.D(\input_filter[0][4] [7]), .CK(n_57_2), 
      .Q(\buffer[6][0][4] [7]), .QN());
   DFF_X1 \buffer_reg[6][0][4][6]  (.D(\input_filter[0][4] [6]), .CK(n_57_2), 
      .Q(\buffer[6][0][4] [6]), .QN());
   DFF_X1 \buffer_reg[6][0][4][5]  (.D(\input_filter[0][4] [5]), .CK(n_57_2), 
      .Q(\buffer[6][0][4] [5]), .QN());
   DFF_X1 \buffer_reg[6][0][4][4]  (.D(\input_filter[0][4] [4]), .CK(n_57_2), 
      .Q(\buffer[6][0][4] [4]), .QN());
   DFF_X1 \buffer_reg[6][0][4][3]  (.D(\input_filter[0][4] [3]), .CK(n_57_2), 
      .Q(\buffer[6][0][4] [3]), .QN());
   DFF_X1 \buffer_reg[6][0][4][2]  (.D(\input_filter[0][4] [2]), .CK(n_57_2), 
      .Q(\buffer[6][0][4] [2]), .QN());
   DFF_X1 \buffer_reg[6][0][4][1]  (.D(\input_filter[0][4] [1]), .CK(n_57_2), 
      .Q(\buffer[6][0][4] [1]), .QN());
   DFF_X1 \buffer_reg[6][0][4][0]  (.D(\input_filter[0][4] [0]), .CK(n_57_2), 
      .Q(\buffer[6][0][4] [0]), .QN());
   CLKGATETST_X1 \clk_gate_buffer_reg[5][0][4]_reg  (.CK(read), .E(n_5), 
      .SE(1'b0), .GCK(n_57_3));
   DFF_X1 \buffer_reg[5][0][4][15]  (.D(\input_filter[0][4] [15]), .CK(n_57_3), 
      .Q(\buffer[5][0][4] [15]), .QN());
   DFF_X1 \buffer_reg[5][0][4][14]  (.D(\input_filter[0][4] [14]), .CK(n_57_3), 
      .Q(\buffer[5][0][4] [14]), .QN());
   DFF_X1 \buffer_reg[5][0][4][13]  (.D(\input_filter[0][4] [13]), .CK(n_57_3), 
      .Q(\buffer[5][0][4] [13]), .QN());
   DFF_X1 \buffer_reg[5][0][4][12]  (.D(\input_filter[0][4] [12]), .CK(n_57_3), 
      .Q(\buffer[5][0][4] [12]), .QN());
   DFF_X1 \buffer_reg[5][0][4][11]  (.D(\input_filter[0][4] [11]), .CK(n_57_3), 
      .Q(\buffer[5][0][4] [11]), .QN());
   DFF_X1 \buffer_reg[5][0][4][10]  (.D(\input_filter[0][4] [10]), .CK(n_57_3), 
      .Q(\buffer[5][0][4] [10]), .QN());
   DFF_X1 \buffer_reg[5][0][4][9]  (.D(\input_filter[0][4] [9]), .CK(n_57_3), 
      .Q(\buffer[5][0][4] [9]), .QN());
   DFF_X1 \buffer_reg[5][0][4][8]  (.D(\input_filter[0][4] [8]), .CK(n_57_3), 
      .Q(\buffer[5][0][4] [8]), .QN());
   DFF_X1 \buffer_reg[5][0][4][7]  (.D(\input_filter[0][4] [7]), .CK(n_57_3), 
      .Q(\buffer[5][0][4] [7]), .QN());
   DFF_X1 \buffer_reg[5][0][4][6]  (.D(\input_filter[0][4] [6]), .CK(n_57_3), 
      .Q(\buffer[5][0][4] [6]), .QN());
   DFF_X1 \buffer_reg[5][0][4][5]  (.D(\input_filter[0][4] [5]), .CK(n_57_3), 
      .Q(\buffer[5][0][4] [5]), .QN());
   DFF_X1 \buffer_reg[5][0][4][4]  (.D(\input_filter[0][4] [4]), .CK(n_57_3), 
      .Q(\buffer[5][0][4] [4]), .QN());
   DFF_X1 \buffer_reg[5][0][4][3]  (.D(\input_filter[0][4] [3]), .CK(n_57_3), 
      .Q(\buffer[5][0][4] [3]), .QN());
   DFF_X1 \buffer_reg[5][0][4][2]  (.D(\input_filter[0][4] [2]), .CK(n_57_3), 
      .Q(\buffer[5][0][4] [2]), .QN());
   DFF_X1 \buffer_reg[5][0][4][1]  (.D(\input_filter[0][4] [1]), .CK(n_57_3), 
      .Q(\buffer[5][0][4] [1]), .QN());
   DFF_X1 \buffer_reg[5][0][4][0]  (.D(\input_filter[0][4] [0]), .CK(n_57_3), 
      .Q(\buffer[5][0][4] [0]), .QN());
   CLKGATETST_X1 \clk_gate_buffer_reg[0][1][2]_reg  (.CK(read), .E(n_0), 
      .SE(1'b0), .GCK(n_57_4));
   CLKGATETST_X1 \clk_gate_buffer_reg[9][1][2]_reg  (.CK(read), .E(n_9), 
      .SE(1'b0), .GCK(n_57_5));
   CLKGATETST_X1 \clk_gate_buffer_reg[10][1][2]_reg  (.CK(read), .E(n_10), 
      .SE(1'b0), .GCK(n_57_6));
   CLKGATETST_X1 \clk_gate_buffer_reg[11][1][2]_reg  (.CK(read), .E(n_11), 
      .SE(1'b0), .GCK(n_57_7));
   CLKGATETST_X1 \clk_gate_buffer_reg[12][1][2]_reg  (.CK(read), .E(n_12), 
      .SE(1'b0), .GCK(n_57_12));
   CLKGATETST_X1 \clk_gate_buffer_reg[13][1][2]_reg  (.CK(read), .E(n_13), 
      .SE(1'b0), .GCK(n_57_13));
   CLKGATETST_X1 \clk_gate_buffer_reg[14][1][2]_reg  (.CK(read), .E(n_14), 
      .SE(1'b0), .GCK(n_57_14));
   CLKGATETST_X1 \clk_gate_buffer_reg[15][1][2]_reg  (.CK(read), .E(n_15), 
      .SE(1'b0), .GCK(n_57_15));
   DFF_X1 \buffer_reg[0][1][3][15]  (.D(\input_filter[1][3] [15]), .CK(n_58_0), 
      .Q(\buffer[0][1][3] [15]), .QN());
   DFF_X1 \buffer_reg[0][1][3][14]  (.D(\input_filter[1][3] [14]), .CK(n_58_0), 
      .Q(\buffer[0][1][3] [14]), .QN());
   DFF_X1 \buffer_reg[0][1][3][13]  (.D(\input_filter[1][3] [13]), .CK(n_58_0), 
      .Q(\buffer[0][1][3] [13]), .QN());
   DFF_X1 \buffer_reg[0][1][3][12]  (.D(\input_filter[1][3] [12]), .CK(n_58_0), 
      .Q(\buffer[0][1][3] [12]), .QN());
   DFF_X1 \buffer_reg[0][1][3][11]  (.D(\input_filter[1][3] [11]), .CK(n_58_0), 
      .Q(\buffer[0][1][3] [11]), .QN());
   DFF_X1 \buffer_reg[0][1][3][10]  (.D(\input_filter[1][3] [10]), .CK(n_58_0), 
      .Q(\buffer[0][1][3] [10]), .QN());
   DFF_X1 \buffer_reg[0][1][3][9]  (.D(\input_filter[1][3] [9]), .CK(n_58_0), 
      .Q(\buffer[0][1][3] [9]), .QN());
   DFF_X1 \buffer_reg[0][1][3][8]  (.D(\input_filter[1][3] [8]), .CK(n_58_0), 
      .Q(\buffer[0][1][3] [8]), .QN());
   DFF_X1 \buffer_reg[0][1][3][7]  (.D(\input_filter[1][3] [7]), .CK(n_58_0), 
      .Q(\buffer[0][1][3] [7]), .QN());
   DFF_X1 \buffer_reg[0][1][3][6]  (.D(\input_filter[1][3] [6]), .CK(n_58_0), 
      .Q(\buffer[0][1][3] [6]), .QN());
   DFF_X1 \buffer_reg[0][1][3][5]  (.D(\input_filter[1][3] [5]), .CK(n_58_0), 
      .Q(\buffer[0][1][3] [5]), .QN());
   DFF_X1 \buffer_reg[0][1][3][4]  (.D(\input_filter[1][3] [4]), .CK(n_58_0), 
      .Q(\buffer[0][1][3] [4]), .QN());
   DFF_X1 \buffer_reg[0][1][3][3]  (.D(\input_filter[1][3] [3]), .CK(n_58_0), 
      .Q(\buffer[0][1][3] [3]), .QN());
   DFF_X1 \buffer_reg[0][1][3][2]  (.D(\input_filter[1][3] [2]), .CK(n_58_0), 
      .Q(\buffer[0][1][3] [2]), .QN());
   DFF_X1 \buffer_reg[0][1][3][1]  (.D(\input_filter[1][3] [1]), .CK(n_58_0), 
      .Q(\buffer[0][1][3] [1]), .QN());
   DFF_X1 \buffer_reg[0][1][3][0]  (.D(\input_filter[1][3] [0]), .CK(n_58_0), 
      .Q(\buffer[0][1][3] [0]), .QN());
   DFF_X1 \buffer_reg[1][1][3][15]  (.D(\input_filter[1][3] [15]), .CK(n_58_1), 
      .Q(\buffer[1][1][3] [15]), .QN());
   DFF_X1 \buffer_reg[1][1][3][14]  (.D(\input_filter[1][3] [14]), .CK(n_58_1), 
      .Q(\buffer[1][1][3] [14]), .QN());
   DFF_X1 \buffer_reg[1][1][3][13]  (.D(\input_filter[1][3] [13]), .CK(n_58_1), 
      .Q(\buffer[1][1][3] [13]), .QN());
   DFF_X1 \buffer_reg[1][1][3][12]  (.D(\input_filter[1][3] [12]), .CK(n_58_1), 
      .Q(\buffer[1][1][3] [12]), .QN());
   DFF_X1 \buffer_reg[1][1][3][11]  (.D(\input_filter[1][3] [11]), .CK(n_58_1), 
      .Q(\buffer[1][1][3] [11]), .QN());
   DFF_X1 \buffer_reg[1][1][3][10]  (.D(\input_filter[1][3] [10]), .CK(n_58_1), 
      .Q(\buffer[1][1][3] [10]), .QN());
   DFF_X1 \buffer_reg[1][1][3][9]  (.D(\input_filter[1][3] [9]), .CK(n_58_1), 
      .Q(\buffer[1][1][3] [9]), .QN());
   DFF_X1 \buffer_reg[1][1][3][8]  (.D(\input_filter[1][3] [8]), .CK(n_58_1), 
      .Q(\buffer[1][1][3] [8]), .QN());
   DFF_X1 \buffer_reg[1][1][3][7]  (.D(\input_filter[1][3] [7]), .CK(n_58_1), 
      .Q(\buffer[1][1][3] [7]), .QN());
   DFF_X1 \buffer_reg[1][1][3][6]  (.D(\input_filter[1][3] [6]), .CK(n_58_1), 
      .Q(\buffer[1][1][3] [6]), .QN());
   DFF_X1 \buffer_reg[1][1][3][5]  (.D(\input_filter[1][3] [5]), .CK(n_58_1), 
      .Q(\buffer[1][1][3] [5]), .QN());
   DFF_X1 \buffer_reg[1][1][3][4]  (.D(\input_filter[1][3] [4]), .CK(n_58_1), 
      .Q(\buffer[1][1][3] [4]), .QN());
   DFF_X1 \buffer_reg[1][1][3][3]  (.D(\input_filter[1][3] [3]), .CK(n_58_1), 
      .Q(\buffer[1][1][3] [3]), .QN());
   DFF_X1 \buffer_reg[1][1][3][2]  (.D(\input_filter[1][3] [2]), .CK(n_58_1), 
      .Q(\buffer[1][1][3] [2]), .QN());
   DFF_X1 \buffer_reg[1][1][3][1]  (.D(\input_filter[1][3] [1]), .CK(n_58_1), 
      .Q(\buffer[1][1][3] [1]), .QN());
   DFF_X1 \buffer_reg[1][1][3][0]  (.D(\input_filter[1][3] [0]), .CK(n_58_1), 
      .Q(\buffer[1][1][3] [0]), .QN());
   DFF_X1 \buffer_reg[2][1][3][15]  (.D(\input_filter[1][3] [15]), .CK(n_58_2), 
      .Q(\buffer[2][1][3] [15]), .QN());
   DFF_X1 \buffer_reg[2][1][3][14]  (.D(\input_filter[1][3] [14]), .CK(n_58_2), 
      .Q(\buffer[2][1][3] [14]), .QN());
   DFF_X1 \buffer_reg[2][1][3][13]  (.D(\input_filter[1][3] [13]), .CK(n_58_2), 
      .Q(\buffer[2][1][3] [13]), .QN());
   DFF_X1 \buffer_reg[2][1][3][12]  (.D(\input_filter[1][3] [12]), .CK(n_58_2), 
      .Q(\buffer[2][1][3] [12]), .QN());
   DFF_X1 \buffer_reg[2][1][3][11]  (.D(\input_filter[1][3] [11]), .CK(n_58_2), 
      .Q(\buffer[2][1][3] [11]), .QN());
   DFF_X1 \buffer_reg[2][1][3][10]  (.D(\input_filter[1][3] [10]), .CK(n_58_2), 
      .Q(\buffer[2][1][3] [10]), .QN());
   DFF_X1 \buffer_reg[2][1][3][9]  (.D(\input_filter[1][3] [9]), .CK(n_58_2), 
      .Q(\buffer[2][1][3] [9]), .QN());
   DFF_X1 \buffer_reg[2][1][3][8]  (.D(\input_filter[1][3] [8]), .CK(n_58_2), 
      .Q(\buffer[2][1][3] [8]), .QN());
   DFF_X1 \buffer_reg[2][1][3][7]  (.D(\input_filter[1][3] [7]), .CK(n_58_2), 
      .Q(\buffer[2][1][3] [7]), .QN());
   DFF_X1 \buffer_reg[2][1][3][6]  (.D(\input_filter[1][3] [6]), .CK(n_58_2), 
      .Q(\buffer[2][1][3] [6]), .QN());
   DFF_X1 \buffer_reg[2][1][3][5]  (.D(\input_filter[1][3] [5]), .CK(n_58_2), 
      .Q(\buffer[2][1][3] [5]), .QN());
   DFF_X1 \buffer_reg[2][1][3][4]  (.D(\input_filter[1][3] [4]), .CK(n_58_2), 
      .Q(\buffer[2][1][3] [4]), .QN());
   DFF_X1 \buffer_reg[2][1][3][3]  (.D(\input_filter[1][3] [3]), .CK(n_58_2), 
      .Q(\buffer[2][1][3] [3]), .QN());
   DFF_X1 \buffer_reg[2][1][3][2]  (.D(\input_filter[1][3] [2]), .CK(n_58_2), 
      .Q(\buffer[2][1][3] [2]), .QN());
   DFF_X1 \buffer_reg[2][1][3][1]  (.D(\input_filter[1][3] [1]), .CK(n_58_2), 
      .Q(\buffer[2][1][3] [1]), .QN());
   DFF_X1 \buffer_reg[2][1][3][0]  (.D(\input_filter[1][3] [0]), .CK(n_58_2), 
      .Q(\buffer[2][1][3] [0]), .QN());
   DFF_X1 \buffer_reg[3][1][3][15]  (.D(\input_filter[1][3] [15]), .CK(n_58_3), 
      .Q(\buffer[3][1][3] [15]), .QN());
   DFF_X1 \buffer_reg[3][1][3][14]  (.D(\input_filter[1][3] [14]), .CK(n_58_3), 
      .Q(\buffer[3][1][3] [14]), .QN());
   DFF_X1 \buffer_reg[3][1][3][13]  (.D(\input_filter[1][3] [13]), .CK(n_58_3), 
      .Q(\buffer[3][1][3] [13]), .QN());
   DFF_X1 \buffer_reg[3][1][3][12]  (.D(\input_filter[1][3] [12]), .CK(n_58_3), 
      .Q(\buffer[3][1][3] [12]), .QN());
   DFF_X1 \buffer_reg[3][1][3][11]  (.D(\input_filter[1][3] [11]), .CK(n_58_3), 
      .Q(\buffer[3][1][3] [11]), .QN());
   DFF_X1 \buffer_reg[3][1][3][10]  (.D(\input_filter[1][3] [10]), .CK(n_58_3), 
      .Q(\buffer[3][1][3] [10]), .QN());
   DFF_X1 \buffer_reg[3][1][3][9]  (.D(\input_filter[1][3] [9]), .CK(n_58_3), 
      .Q(\buffer[3][1][3] [9]), .QN());
   DFF_X1 \buffer_reg[3][1][3][8]  (.D(\input_filter[1][3] [8]), .CK(n_58_3), 
      .Q(\buffer[3][1][3] [8]), .QN());
   DFF_X1 \buffer_reg[3][1][3][7]  (.D(\input_filter[1][3] [7]), .CK(n_58_3), 
      .Q(\buffer[3][1][3] [7]), .QN());
   DFF_X1 \buffer_reg[3][1][3][6]  (.D(\input_filter[1][3] [6]), .CK(n_58_3), 
      .Q(\buffer[3][1][3] [6]), .QN());
   DFF_X1 \buffer_reg[3][1][3][5]  (.D(\input_filter[1][3] [5]), .CK(n_58_3), 
      .Q(\buffer[3][1][3] [5]), .QN());
   DFF_X1 \buffer_reg[3][1][3][4]  (.D(\input_filter[1][3] [4]), .CK(n_58_3), 
      .Q(\buffer[3][1][3] [4]), .QN());
   DFF_X1 \buffer_reg[3][1][3][3]  (.D(\input_filter[1][3] [3]), .CK(n_58_3), 
      .Q(\buffer[3][1][3] [3]), .QN());
   DFF_X1 \buffer_reg[3][1][3][2]  (.D(\input_filter[1][3] [2]), .CK(n_58_3), 
      .Q(\buffer[3][1][3] [2]), .QN());
   DFF_X1 \buffer_reg[3][1][3][1]  (.D(\input_filter[1][3] [1]), .CK(n_58_3), 
      .Q(\buffer[3][1][3] [1]), .QN());
   DFF_X1 \buffer_reg[3][1][3][0]  (.D(\input_filter[1][3] [0]), .CK(n_58_3), 
      .Q(\buffer[3][1][3] [0]), .QN());
   DFF_X1 \buffer_reg[4][1][3][15]  (.D(\input_filter[1][3] [15]), .CK(n_58_4), 
      .Q(\buffer[4][1][3] [15]), .QN());
   DFF_X1 \buffer_reg[4][1][3][14]  (.D(\input_filter[1][3] [14]), .CK(n_58_4), 
      .Q(\buffer[4][1][3] [14]), .QN());
   DFF_X1 \buffer_reg[4][1][3][13]  (.D(\input_filter[1][3] [13]), .CK(n_58_4), 
      .Q(\buffer[4][1][3] [13]), .QN());
   DFF_X1 \buffer_reg[4][1][3][12]  (.D(\input_filter[1][3] [12]), .CK(n_58_4), 
      .Q(\buffer[4][1][3] [12]), .QN());
   DFF_X1 \buffer_reg[4][1][3][11]  (.D(\input_filter[1][3] [11]), .CK(n_58_4), 
      .Q(\buffer[4][1][3] [11]), .QN());
   DFF_X1 \buffer_reg[4][1][3][10]  (.D(\input_filter[1][3] [10]), .CK(n_58_4), 
      .Q(\buffer[4][1][3] [10]), .QN());
   DFF_X1 \buffer_reg[4][1][3][9]  (.D(\input_filter[1][3] [9]), .CK(n_58_4), 
      .Q(\buffer[4][1][3] [9]), .QN());
   DFF_X1 \buffer_reg[4][1][3][8]  (.D(\input_filter[1][3] [8]), .CK(n_58_4), 
      .Q(\buffer[4][1][3] [8]), .QN());
   DFF_X1 \buffer_reg[4][1][3][7]  (.D(\input_filter[1][3] [7]), .CK(n_58_4), 
      .Q(\buffer[4][1][3] [7]), .QN());
   DFF_X1 \buffer_reg[4][1][3][6]  (.D(\input_filter[1][3] [6]), .CK(n_58_4), 
      .Q(\buffer[4][1][3] [6]), .QN());
   DFF_X1 \buffer_reg[4][1][3][5]  (.D(\input_filter[1][3] [5]), .CK(n_58_4), 
      .Q(\buffer[4][1][3] [5]), .QN());
   DFF_X1 \buffer_reg[4][1][3][4]  (.D(\input_filter[1][3] [4]), .CK(n_58_4), 
      .Q(\buffer[4][1][3] [4]), .QN());
   DFF_X1 \buffer_reg[4][1][3][3]  (.D(\input_filter[1][3] [3]), .CK(n_58_4), 
      .Q(\buffer[4][1][3] [3]), .QN());
   DFF_X1 \buffer_reg[4][1][3][2]  (.D(\input_filter[1][3] [2]), .CK(n_58_4), 
      .Q(\buffer[4][1][3] [2]), .QN());
   DFF_X1 \buffer_reg[4][1][3][1]  (.D(\input_filter[1][3] [1]), .CK(n_58_4), 
      .Q(\buffer[4][1][3] [1]), .QN());
   DFF_X1 \buffer_reg[4][1][3][0]  (.D(\input_filter[1][3] [0]), .CK(n_58_4), 
      .Q(\buffer[4][1][3] [0]), .QN());
   DFF_X1 \buffer_reg[5][1][3][15]  (.D(\input_filter[1][3] [15]), .CK(n_58_5), 
      .Q(\buffer[5][1][3] [15]), .QN());
   DFF_X1 \buffer_reg[5][1][3][14]  (.D(\input_filter[1][3] [14]), .CK(n_58_5), 
      .Q(\buffer[5][1][3] [14]), .QN());
   DFF_X1 \buffer_reg[5][1][3][13]  (.D(\input_filter[1][3] [13]), .CK(n_58_5), 
      .Q(\buffer[5][1][3] [13]), .QN());
   DFF_X1 \buffer_reg[5][1][3][12]  (.D(\input_filter[1][3] [12]), .CK(n_58_5), 
      .Q(\buffer[5][1][3] [12]), .QN());
   DFF_X1 \buffer_reg[5][1][3][11]  (.D(\input_filter[1][3] [11]), .CK(n_58_5), 
      .Q(\buffer[5][1][3] [11]), .QN());
   DFF_X1 \buffer_reg[5][1][3][10]  (.D(\input_filter[1][3] [10]), .CK(n_58_5), 
      .Q(\buffer[5][1][3] [10]), .QN());
   DFF_X1 \buffer_reg[5][1][3][9]  (.D(\input_filter[1][3] [9]), .CK(n_58_5), 
      .Q(\buffer[5][1][3] [9]), .QN());
   DFF_X1 \buffer_reg[5][1][3][8]  (.D(\input_filter[1][3] [8]), .CK(n_58_5), 
      .Q(\buffer[5][1][3] [8]), .QN());
   DFF_X1 \buffer_reg[5][1][3][7]  (.D(\input_filter[1][3] [7]), .CK(n_58_5), 
      .Q(\buffer[5][1][3] [7]), .QN());
   DFF_X1 \buffer_reg[5][1][3][6]  (.D(\input_filter[1][3] [6]), .CK(n_58_5), 
      .Q(\buffer[5][1][3] [6]), .QN());
   DFF_X1 \buffer_reg[5][1][3][5]  (.D(\input_filter[1][3] [5]), .CK(n_58_5), 
      .Q(\buffer[5][1][3] [5]), .QN());
   DFF_X1 \buffer_reg[5][1][3][4]  (.D(\input_filter[1][3] [4]), .CK(n_58_5), 
      .Q(\buffer[5][1][3] [4]), .QN());
   DFF_X1 \buffer_reg[5][1][3][3]  (.D(\input_filter[1][3] [3]), .CK(n_58_5), 
      .Q(\buffer[5][1][3] [3]), .QN());
   DFF_X1 \buffer_reg[5][1][3][2]  (.D(\input_filter[1][3] [2]), .CK(n_58_5), 
      .Q(\buffer[5][1][3] [2]), .QN());
   DFF_X1 \buffer_reg[5][1][3][1]  (.D(\input_filter[1][3] [1]), .CK(n_58_5), 
      .Q(\buffer[5][1][3] [1]), .QN());
   DFF_X1 \buffer_reg[5][1][3][0]  (.D(\input_filter[1][3] [0]), .CK(n_58_5), 
      .Q(\buffer[5][1][3] [0]), .QN());
   CLKGATETST_X1 \clk_gate_buffer_reg[6][1][3]_reg  (.CK(read), .E(n_6), 
      .SE(1'b0), .GCK(n_58_6));
   DFF_X1 \buffer_reg[6][1][3][15]  (.D(\input_filter[1][3] [15]), .CK(n_58_6), 
      .Q(\buffer[6][1][3] [15]), .QN());
   DFF_X1 \buffer_reg[6][1][3][14]  (.D(\input_filter[1][3] [14]), .CK(n_58_6), 
      .Q(\buffer[6][1][3] [14]), .QN());
   DFF_X1 \buffer_reg[6][1][3][13]  (.D(\input_filter[1][3] [13]), .CK(n_58_6), 
      .Q(\buffer[6][1][3] [13]), .QN());
   DFF_X1 \buffer_reg[6][1][3][12]  (.D(\input_filter[1][3] [12]), .CK(n_58_6), 
      .Q(\buffer[6][1][3] [12]), .QN());
   DFF_X1 \buffer_reg[6][1][3][11]  (.D(\input_filter[1][3] [11]), .CK(n_58_6), 
      .Q(\buffer[6][1][3] [11]), .QN());
   DFF_X1 \buffer_reg[6][1][3][10]  (.D(\input_filter[1][3] [10]), .CK(n_58_6), 
      .Q(\buffer[6][1][3] [10]), .QN());
   DFF_X1 \buffer_reg[6][1][3][9]  (.D(\input_filter[1][3] [9]), .CK(n_58_6), 
      .Q(\buffer[6][1][3] [9]), .QN());
   DFF_X1 \buffer_reg[6][1][3][8]  (.D(\input_filter[1][3] [8]), .CK(n_58_6), 
      .Q(\buffer[6][1][3] [8]), .QN());
   DFF_X1 \buffer_reg[6][1][3][7]  (.D(\input_filter[1][3] [7]), .CK(n_58_6), 
      .Q(\buffer[6][1][3] [7]), .QN());
   DFF_X1 \buffer_reg[6][1][3][6]  (.D(\input_filter[1][3] [6]), .CK(n_58_6), 
      .Q(\buffer[6][1][3] [6]), .QN());
   DFF_X1 \buffer_reg[6][1][3][5]  (.D(\input_filter[1][3] [5]), .CK(n_58_6), 
      .Q(\buffer[6][1][3] [5]), .QN());
   DFF_X1 \buffer_reg[6][1][3][4]  (.D(\input_filter[1][3] [4]), .CK(n_58_6), 
      .Q(\buffer[6][1][3] [4]), .QN());
   DFF_X1 \buffer_reg[6][1][3][3]  (.D(\input_filter[1][3] [3]), .CK(n_58_6), 
      .Q(\buffer[6][1][3] [3]), .QN());
   DFF_X1 \buffer_reg[6][1][3][2]  (.D(\input_filter[1][3] [2]), .CK(n_58_6), 
      .Q(\buffer[6][1][3] [2]), .QN());
   DFF_X1 \buffer_reg[6][1][3][1]  (.D(\input_filter[1][3] [1]), .CK(n_58_6), 
      .Q(\buffer[6][1][3] [1]), .QN());
   DFF_X1 \buffer_reg[6][1][3][0]  (.D(\input_filter[1][3] [0]), .CK(n_58_6), 
      .Q(\buffer[6][1][3] [0]), .QN());
   DFF_X1 \buffer_reg[7][1][3][15]  (.D(\input_filter[1][3] [15]), .CK(n_58_7), 
      .Q(\buffer[7][1][3] [15]), .QN());
   DFF_X1 \buffer_reg[7][1][3][14]  (.D(\input_filter[1][3] [14]), .CK(n_58_7), 
      .Q(\buffer[7][1][3] [14]), .QN());
   DFF_X1 \buffer_reg[7][1][3][13]  (.D(\input_filter[1][3] [13]), .CK(n_58_7), 
      .Q(\buffer[7][1][3] [13]), .QN());
   DFF_X1 \buffer_reg[7][1][3][12]  (.D(\input_filter[1][3] [12]), .CK(n_58_7), 
      .Q(\buffer[7][1][3] [12]), .QN());
   DFF_X1 \buffer_reg[7][1][3][11]  (.D(\input_filter[1][3] [11]), .CK(n_58_7), 
      .Q(\buffer[7][1][3] [11]), .QN());
   DFF_X1 \buffer_reg[7][1][3][10]  (.D(\input_filter[1][3] [10]), .CK(n_58_7), 
      .Q(\buffer[7][1][3] [10]), .QN());
   DFF_X1 \buffer_reg[7][1][3][9]  (.D(\input_filter[1][3] [9]), .CK(n_58_7), 
      .Q(\buffer[7][1][3] [9]), .QN());
   DFF_X1 \buffer_reg[7][1][3][8]  (.D(\input_filter[1][3] [8]), .CK(n_58_7), 
      .Q(\buffer[7][1][3] [8]), .QN());
   DFF_X1 \buffer_reg[7][1][3][7]  (.D(\input_filter[1][3] [7]), .CK(n_58_7), 
      .Q(\buffer[7][1][3] [7]), .QN());
   DFF_X1 \buffer_reg[7][1][3][6]  (.D(\input_filter[1][3] [6]), .CK(n_58_7), 
      .Q(\buffer[7][1][3] [6]), .QN());
   DFF_X1 \buffer_reg[7][1][3][5]  (.D(\input_filter[1][3] [5]), .CK(n_58_7), 
      .Q(\buffer[7][1][3] [5]), .QN());
   DFF_X1 \buffer_reg[7][1][3][4]  (.D(\input_filter[1][3] [4]), .CK(n_58_7), 
      .Q(\buffer[7][1][3] [4]), .QN());
   DFF_X1 \buffer_reg[7][1][3][3]  (.D(\input_filter[1][3] [3]), .CK(n_58_7), 
      .Q(\buffer[7][1][3] [3]), .QN());
   DFF_X1 \buffer_reg[7][1][3][2]  (.D(\input_filter[1][3] [2]), .CK(n_58_7), 
      .Q(\buffer[7][1][3] [2]), .QN());
   DFF_X1 \buffer_reg[7][1][3][1]  (.D(\input_filter[1][3] [1]), .CK(n_58_7), 
      .Q(\buffer[7][1][3] [1]), .QN());
   DFF_X1 \buffer_reg[7][1][3][0]  (.D(\input_filter[1][3] [0]), .CK(n_58_7), 
      .Q(\buffer[7][1][3] [0]), .QN());
   DFF_X1 \buffer_reg[8][1][3][15]  (.D(\input_filter[1][3] [15]), .CK(n_58_8), 
      .Q(\buffer[8][1][3] [15]), .QN());
   DFF_X1 \buffer_reg[8][1][3][14]  (.D(\input_filter[1][3] [14]), .CK(n_58_8), 
      .Q(\buffer[8][1][3] [14]), .QN());
   DFF_X1 \buffer_reg[8][1][3][13]  (.D(\input_filter[1][3] [13]), .CK(n_58_8), 
      .Q(\buffer[8][1][3] [13]), .QN());
   DFF_X1 \buffer_reg[8][1][3][12]  (.D(\input_filter[1][3] [12]), .CK(n_58_8), 
      .Q(\buffer[8][1][3] [12]), .QN());
   DFF_X1 \buffer_reg[8][1][3][11]  (.D(\input_filter[1][3] [11]), .CK(n_58_8), 
      .Q(\buffer[8][1][3] [11]), .QN());
   DFF_X1 \buffer_reg[8][1][3][10]  (.D(\input_filter[1][3] [10]), .CK(n_58_8), 
      .Q(\buffer[8][1][3] [10]), .QN());
   DFF_X1 \buffer_reg[8][1][3][9]  (.D(\input_filter[1][3] [9]), .CK(n_58_8), 
      .Q(\buffer[8][1][3] [9]), .QN());
   DFF_X1 \buffer_reg[8][1][3][8]  (.D(\input_filter[1][3] [8]), .CK(n_58_8), 
      .Q(\buffer[8][1][3] [8]), .QN());
   DFF_X1 \buffer_reg[8][1][3][7]  (.D(\input_filter[1][3] [7]), .CK(n_58_8), 
      .Q(\buffer[8][1][3] [7]), .QN());
   DFF_X1 \buffer_reg[8][1][3][6]  (.D(\input_filter[1][3] [6]), .CK(n_58_8), 
      .Q(\buffer[8][1][3] [6]), .QN());
   DFF_X1 \buffer_reg[8][1][3][5]  (.D(\input_filter[1][3] [5]), .CK(n_58_8), 
      .Q(\buffer[8][1][3] [5]), .QN());
   DFF_X1 \buffer_reg[8][1][3][4]  (.D(\input_filter[1][3] [4]), .CK(n_58_8), 
      .Q(\buffer[8][1][3] [4]), .QN());
   DFF_X1 \buffer_reg[8][1][3][3]  (.D(\input_filter[1][3] [3]), .CK(n_58_8), 
      .Q(\buffer[8][1][3] [3]), .QN());
   DFF_X1 \buffer_reg[8][1][3][2]  (.D(\input_filter[1][3] [2]), .CK(n_58_8), 
      .Q(\buffer[8][1][3] [2]), .QN());
   DFF_X1 \buffer_reg[8][1][3][1]  (.D(\input_filter[1][3] [1]), .CK(n_58_8), 
      .Q(\buffer[8][1][3] [1]), .QN());
   DFF_X1 \buffer_reg[8][1][3][0]  (.D(\input_filter[1][3] [0]), .CK(n_58_8), 
      .Q(\buffer[8][1][3] [0]), .QN());
   DFF_X1 \buffer_reg[9][1][3][15]  (.D(\input_filter[1][3] [15]), .CK(n_58_9), 
      .Q(\buffer[9][1][3] [15]), .QN());
   DFF_X1 \buffer_reg[9][1][3][14]  (.D(\input_filter[1][3] [14]), .CK(n_58_9), 
      .Q(\buffer[9][1][3] [14]), .QN());
   DFF_X1 \buffer_reg[9][1][3][13]  (.D(\input_filter[1][3] [13]), .CK(n_58_9), 
      .Q(\buffer[9][1][3] [13]), .QN());
   DFF_X1 \buffer_reg[9][1][3][12]  (.D(\input_filter[1][3] [12]), .CK(n_58_9), 
      .Q(\buffer[9][1][3] [12]), .QN());
   DFF_X1 \buffer_reg[9][1][3][11]  (.D(\input_filter[1][3] [11]), .CK(n_58_9), 
      .Q(\buffer[9][1][3] [11]), .QN());
   DFF_X1 \buffer_reg[9][1][3][10]  (.D(\input_filter[1][3] [10]), .CK(n_58_9), 
      .Q(\buffer[9][1][3] [10]), .QN());
   DFF_X1 \buffer_reg[9][1][3][9]  (.D(\input_filter[1][3] [9]), .CK(n_58_9), 
      .Q(\buffer[9][1][3] [9]), .QN());
   DFF_X1 \buffer_reg[9][1][3][8]  (.D(\input_filter[1][3] [8]), .CK(n_58_9), 
      .Q(\buffer[9][1][3] [8]), .QN());
   DFF_X1 \buffer_reg[9][1][3][7]  (.D(\input_filter[1][3] [7]), .CK(n_58_9), 
      .Q(\buffer[9][1][3] [7]), .QN());
   DFF_X1 \buffer_reg[9][1][3][6]  (.D(\input_filter[1][3] [6]), .CK(n_58_9), 
      .Q(\buffer[9][1][3] [6]), .QN());
   DFF_X1 \buffer_reg[9][1][3][5]  (.D(\input_filter[1][3] [5]), .CK(n_58_9), 
      .Q(\buffer[9][1][3] [5]), .QN());
   DFF_X1 \buffer_reg[9][1][3][4]  (.D(\input_filter[1][3] [4]), .CK(n_58_9), 
      .Q(\buffer[9][1][3] [4]), .QN());
   DFF_X1 \buffer_reg[9][1][3][3]  (.D(\input_filter[1][3] [3]), .CK(n_58_9), 
      .Q(\buffer[9][1][3] [3]), .QN());
   DFF_X1 \buffer_reg[9][1][3][2]  (.D(\input_filter[1][3] [2]), .CK(n_58_9), 
      .Q(\buffer[9][1][3] [2]), .QN());
   DFF_X1 \buffer_reg[9][1][3][1]  (.D(\input_filter[1][3] [1]), .CK(n_58_9), 
      .Q(\buffer[9][1][3] [1]), .QN());
   DFF_X1 \buffer_reg[9][1][3][0]  (.D(\input_filter[1][3] [0]), .CK(n_58_9), 
      .Q(\buffer[9][1][3] [0]), .QN());
   DFF_X1 \buffer_reg[10][1][3][15]  (.D(\input_filter[1][3] [15]), .CK(n_58_10), 
      .Q(\buffer[10][1][3] [15]), .QN());
   DFF_X1 \buffer_reg[10][1][3][14]  (.D(\input_filter[1][3] [14]), .CK(n_58_10), 
      .Q(\buffer[10][1][3] [14]), .QN());
   DFF_X1 \buffer_reg[10][1][3][13]  (.D(\input_filter[1][3] [13]), .CK(n_58_10), 
      .Q(\buffer[10][1][3] [13]), .QN());
   DFF_X1 \buffer_reg[10][1][3][12]  (.D(\input_filter[1][3] [12]), .CK(n_58_10), 
      .Q(\buffer[10][1][3] [12]), .QN());
   DFF_X1 \buffer_reg[10][1][3][11]  (.D(\input_filter[1][3] [11]), .CK(n_58_10), 
      .Q(\buffer[10][1][3] [11]), .QN());
   DFF_X1 \buffer_reg[10][1][3][10]  (.D(\input_filter[1][3] [10]), .CK(n_58_10), 
      .Q(\buffer[10][1][3] [10]), .QN());
   DFF_X1 \buffer_reg[10][1][3][9]  (.D(\input_filter[1][3] [9]), .CK(n_58_10), 
      .Q(\buffer[10][1][3] [9]), .QN());
   DFF_X1 \buffer_reg[10][1][3][8]  (.D(\input_filter[1][3] [8]), .CK(n_58_10), 
      .Q(\buffer[10][1][3] [8]), .QN());
   DFF_X1 \buffer_reg[10][1][3][7]  (.D(\input_filter[1][3] [7]), .CK(n_58_10), 
      .Q(\buffer[10][1][3] [7]), .QN());
   DFF_X1 \buffer_reg[10][1][3][6]  (.D(\input_filter[1][3] [6]), .CK(n_58_10), 
      .Q(\buffer[10][1][3] [6]), .QN());
   DFF_X1 \buffer_reg[10][1][3][5]  (.D(\input_filter[1][3] [5]), .CK(n_58_10), 
      .Q(\buffer[10][1][3] [5]), .QN());
   DFF_X1 \buffer_reg[10][1][3][4]  (.D(\input_filter[1][3] [4]), .CK(n_58_10), 
      .Q(\buffer[10][1][3] [4]), .QN());
   DFF_X1 \buffer_reg[10][1][3][3]  (.D(\input_filter[1][3] [3]), .CK(n_58_10), 
      .Q(\buffer[10][1][3] [3]), .QN());
   DFF_X1 \buffer_reg[10][1][3][2]  (.D(\input_filter[1][3] [2]), .CK(n_58_10), 
      .Q(\buffer[10][1][3] [2]), .QN());
   DFF_X1 \buffer_reg[10][1][3][1]  (.D(\input_filter[1][3] [1]), .CK(n_58_10), 
      .Q(\buffer[10][1][3] [1]), .QN());
   DFF_X1 \buffer_reg[10][1][3][0]  (.D(\input_filter[1][3] [0]), .CK(n_58_10), 
      .Q(\buffer[10][1][3] [0]), .QN());
   DFF_X1 \buffer_reg[11][1][3][15]  (.D(\input_filter[1][3] [15]), .CK(n_58_11), 
      .Q(\buffer[11][1][3] [15]), .QN());
   DFF_X1 \buffer_reg[11][1][3][14]  (.D(\input_filter[1][3] [14]), .CK(n_58_11), 
      .Q(\buffer[11][1][3] [14]), .QN());
   DFF_X1 \buffer_reg[11][1][3][13]  (.D(\input_filter[1][3] [13]), .CK(n_58_11), 
      .Q(\buffer[11][1][3] [13]), .QN());
   DFF_X1 \buffer_reg[11][1][3][12]  (.D(\input_filter[1][3] [12]), .CK(n_58_11), 
      .Q(\buffer[11][1][3] [12]), .QN());
   DFF_X1 \buffer_reg[11][1][3][11]  (.D(\input_filter[1][3] [11]), .CK(n_58_11), 
      .Q(\buffer[11][1][3] [11]), .QN());
   DFF_X1 \buffer_reg[11][1][3][10]  (.D(\input_filter[1][3] [10]), .CK(n_58_11), 
      .Q(\buffer[11][1][3] [10]), .QN());
   DFF_X1 \buffer_reg[11][1][3][9]  (.D(\input_filter[1][3] [9]), .CK(n_58_11), 
      .Q(\buffer[11][1][3] [9]), .QN());
   DFF_X1 \buffer_reg[11][1][3][8]  (.D(\input_filter[1][3] [8]), .CK(n_58_11), 
      .Q(\buffer[11][1][3] [8]), .QN());
   DFF_X1 \buffer_reg[11][1][3][7]  (.D(\input_filter[1][3] [7]), .CK(n_58_11), 
      .Q(\buffer[11][1][3] [7]), .QN());
   DFF_X1 \buffer_reg[11][1][3][6]  (.D(\input_filter[1][3] [6]), .CK(n_58_11), 
      .Q(\buffer[11][1][3] [6]), .QN());
   DFF_X1 \buffer_reg[11][1][3][5]  (.D(\input_filter[1][3] [5]), .CK(n_58_11), 
      .Q(\buffer[11][1][3] [5]), .QN());
   DFF_X1 \buffer_reg[11][1][3][4]  (.D(\input_filter[1][3] [4]), .CK(n_58_11), 
      .Q(\buffer[11][1][3] [4]), .QN());
   DFF_X1 \buffer_reg[11][1][3][3]  (.D(\input_filter[1][3] [3]), .CK(n_58_11), 
      .Q(\buffer[11][1][3] [3]), .QN());
   DFF_X1 \buffer_reg[11][1][3][2]  (.D(\input_filter[1][3] [2]), .CK(n_58_11), 
      .Q(\buffer[11][1][3] [2]), .QN());
   DFF_X1 \buffer_reg[11][1][3][1]  (.D(\input_filter[1][3] [1]), .CK(n_58_11), 
      .Q(\buffer[11][1][3] [1]), .QN());
   DFF_X1 \buffer_reg[11][1][3][0]  (.D(\input_filter[1][3] [0]), .CK(n_58_11), 
      .Q(\buffer[11][1][3] [0]), .QN());
   DFF_X1 \buffer_reg[12][1][3][15]  (.D(\input_filter[1][3] [15]), .CK(n_58_12), 
      .Q(\buffer[12][1][3] [15]), .QN());
   DFF_X1 \buffer_reg[12][1][3][14]  (.D(\input_filter[1][3] [14]), .CK(n_58_12), 
      .Q(\buffer[12][1][3] [14]), .QN());
   DFF_X1 \buffer_reg[12][1][3][13]  (.D(\input_filter[1][3] [13]), .CK(n_58_12), 
      .Q(\buffer[12][1][3] [13]), .QN());
   DFF_X1 \buffer_reg[12][1][3][12]  (.D(\input_filter[1][3] [12]), .CK(n_58_12), 
      .Q(\buffer[12][1][3] [12]), .QN());
   DFF_X1 \buffer_reg[12][1][3][11]  (.D(\input_filter[1][3] [11]), .CK(n_58_12), 
      .Q(\buffer[12][1][3] [11]), .QN());
   DFF_X1 \buffer_reg[12][1][3][10]  (.D(\input_filter[1][3] [10]), .CK(n_58_12), 
      .Q(\buffer[12][1][3] [10]), .QN());
   DFF_X1 \buffer_reg[12][1][3][9]  (.D(\input_filter[1][3] [9]), .CK(n_58_12), 
      .Q(\buffer[12][1][3] [9]), .QN());
   DFF_X1 \buffer_reg[12][1][3][8]  (.D(\input_filter[1][3] [8]), .CK(n_58_12), 
      .Q(\buffer[12][1][3] [8]), .QN());
   DFF_X1 \buffer_reg[12][1][3][7]  (.D(\input_filter[1][3] [7]), .CK(n_58_12), 
      .Q(\buffer[12][1][3] [7]), .QN());
   DFF_X1 \buffer_reg[12][1][3][6]  (.D(\input_filter[1][3] [6]), .CK(n_58_12), 
      .Q(\buffer[12][1][3] [6]), .QN());
   DFF_X1 \buffer_reg[12][1][3][5]  (.D(\input_filter[1][3] [5]), .CK(n_58_12), 
      .Q(\buffer[12][1][3] [5]), .QN());
   DFF_X1 \buffer_reg[12][1][3][4]  (.D(\input_filter[1][3] [4]), .CK(n_58_12), 
      .Q(\buffer[12][1][3] [4]), .QN());
   DFF_X1 \buffer_reg[12][1][3][3]  (.D(\input_filter[1][3] [3]), .CK(n_58_12), 
      .Q(\buffer[12][1][3] [3]), .QN());
   DFF_X1 \buffer_reg[12][1][3][2]  (.D(\input_filter[1][3] [2]), .CK(n_58_12), 
      .Q(\buffer[12][1][3] [2]), .QN());
   DFF_X1 \buffer_reg[12][1][3][1]  (.D(\input_filter[1][3] [1]), .CK(n_58_12), 
      .Q(\buffer[12][1][3] [1]), .QN());
   DFF_X1 \buffer_reg[12][1][3][0]  (.D(\input_filter[1][3] [0]), .CK(n_58_12), 
      .Q(\buffer[12][1][3] [0]), .QN());
   DFF_X1 \buffer_reg[13][1][3][15]  (.D(\input_filter[1][3] [15]), .CK(n_58_13), 
      .Q(\buffer[13][1][3] [15]), .QN());
   DFF_X1 \buffer_reg[13][1][3][14]  (.D(\input_filter[1][3] [14]), .CK(n_58_13), 
      .Q(\buffer[13][1][3] [14]), .QN());
   DFF_X1 \buffer_reg[13][1][3][13]  (.D(\input_filter[1][3] [13]), .CK(n_58_13), 
      .Q(\buffer[13][1][3] [13]), .QN());
   DFF_X1 \buffer_reg[13][1][3][12]  (.D(\input_filter[1][3] [12]), .CK(n_58_13), 
      .Q(\buffer[13][1][3] [12]), .QN());
   DFF_X1 \buffer_reg[13][1][3][11]  (.D(\input_filter[1][3] [11]), .CK(n_58_13), 
      .Q(\buffer[13][1][3] [11]), .QN());
   DFF_X1 \buffer_reg[13][1][3][10]  (.D(\input_filter[1][3] [10]), .CK(n_58_13), 
      .Q(\buffer[13][1][3] [10]), .QN());
   DFF_X1 \buffer_reg[13][1][3][9]  (.D(\input_filter[1][3] [9]), .CK(n_58_13), 
      .Q(\buffer[13][1][3] [9]), .QN());
   DFF_X1 \buffer_reg[13][1][3][8]  (.D(\input_filter[1][3] [8]), .CK(n_58_13), 
      .Q(\buffer[13][1][3] [8]), .QN());
   DFF_X1 \buffer_reg[13][1][3][7]  (.D(\input_filter[1][3] [7]), .CK(n_58_13), 
      .Q(\buffer[13][1][3] [7]), .QN());
   DFF_X1 \buffer_reg[13][1][3][6]  (.D(\input_filter[1][3] [6]), .CK(n_58_13), 
      .Q(\buffer[13][1][3] [6]), .QN());
   DFF_X1 \buffer_reg[13][1][3][5]  (.D(\input_filter[1][3] [5]), .CK(n_58_13), 
      .Q(\buffer[13][1][3] [5]), .QN());
   DFF_X1 \buffer_reg[13][1][3][4]  (.D(\input_filter[1][3] [4]), .CK(n_58_13), 
      .Q(\buffer[13][1][3] [4]), .QN());
   DFF_X1 \buffer_reg[13][1][3][3]  (.D(\input_filter[1][3] [3]), .CK(n_58_13), 
      .Q(\buffer[13][1][3] [3]), .QN());
   DFF_X1 \buffer_reg[13][1][3][2]  (.D(\input_filter[1][3] [2]), .CK(n_58_13), 
      .Q(\buffer[13][1][3] [2]), .QN());
   DFF_X1 \buffer_reg[13][1][3][1]  (.D(\input_filter[1][3] [1]), .CK(n_58_13), 
      .Q(\buffer[13][1][3] [1]), .QN());
   DFF_X1 \buffer_reg[13][1][3][0]  (.D(\input_filter[1][3] [0]), .CK(n_58_13), 
      .Q(\buffer[13][1][3] [0]), .QN());
   DFF_X1 \buffer_reg[14][1][3][15]  (.D(\input_filter[1][3] [15]), .CK(n_58_14), 
      .Q(\buffer[14][1][3] [15]), .QN());
   DFF_X1 \buffer_reg[14][1][3][14]  (.D(\input_filter[1][3] [14]), .CK(n_58_14), 
      .Q(\buffer[14][1][3] [14]), .QN());
   DFF_X1 \buffer_reg[14][1][3][13]  (.D(\input_filter[1][3] [13]), .CK(n_58_14), 
      .Q(\buffer[14][1][3] [13]), .QN());
   DFF_X1 \buffer_reg[14][1][3][12]  (.D(\input_filter[1][3] [12]), .CK(n_58_14), 
      .Q(\buffer[14][1][3] [12]), .QN());
   DFF_X1 \buffer_reg[14][1][3][11]  (.D(\input_filter[1][3] [11]), .CK(n_58_14), 
      .Q(\buffer[14][1][3] [11]), .QN());
   DFF_X1 \buffer_reg[14][1][3][10]  (.D(\input_filter[1][3] [10]), .CK(n_58_14), 
      .Q(\buffer[14][1][3] [10]), .QN());
   DFF_X1 \buffer_reg[14][1][3][9]  (.D(\input_filter[1][3] [9]), .CK(n_58_14), 
      .Q(\buffer[14][1][3] [9]), .QN());
   DFF_X1 \buffer_reg[14][1][3][8]  (.D(\input_filter[1][3] [8]), .CK(n_58_14), 
      .Q(\buffer[14][1][3] [8]), .QN());
   DFF_X1 \buffer_reg[14][1][3][7]  (.D(\input_filter[1][3] [7]), .CK(n_58_14), 
      .Q(\buffer[14][1][3] [7]), .QN());
   DFF_X1 \buffer_reg[14][1][3][6]  (.D(\input_filter[1][3] [6]), .CK(n_58_14), 
      .Q(\buffer[14][1][3] [6]), .QN());
   DFF_X1 \buffer_reg[14][1][3][5]  (.D(\input_filter[1][3] [5]), .CK(n_58_14), 
      .Q(\buffer[14][1][3] [5]), .QN());
   DFF_X1 \buffer_reg[14][1][3][4]  (.D(\input_filter[1][3] [4]), .CK(n_58_14), 
      .Q(\buffer[14][1][3] [4]), .QN());
   DFF_X1 \buffer_reg[14][1][3][3]  (.D(\input_filter[1][3] [3]), .CK(n_58_14), 
      .Q(\buffer[14][1][3] [3]), .QN());
   DFF_X1 \buffer_reg[14][1][3][2]  (.D(\input_filter[1][3] [2]), .CK(n_58_14), 
      .Q(\buffer[14][1][3] [2]), .QN());
   DFF_X1 \buffer_reg[14][1][3][1]  (.D(\input_filter[1][3] [1]), .CK(n_58_14), 
      .Q(\buffer[14][1][3] [1]), .QN());
   DFF_X1 \buffer_reg[14][1][3][0]  (.D(\input_filter[1][3] [0]), .CK(n_58_14), 
      .Q(\buffer[14][1][3] [0]), .QN());
   CLKGATETST_X1 \clk_gate_buffer_reg[15][1][3]_reg  (.CK(read), .E(n_15), 
      .SE(1'b0), .GCK(n_58_15));
   DFF_X1 \buffer_reg[15][1][3][15]  (.D(\input_filter[1][3] [15]), .CK(n_58_15), 
      .Q(\buffer[15][1][3] [15]), .QN());
   DFF_X1 \buffer_reg[15][1][3][14]  (.D(\input_filter[1][3] [14]), .CK(n_58_15), 
      .Q(\buffer[15][1][3] [14]), .QN());
   DFF_X1 \buffer_reg[15][1][3][13]  (.D(\input_filter[1][3] [13]), .CK(n_58_15), 
      .Q(\buffer[15][1][3] [13]), .QN());
   DFF_X1 \buffer_reg[15][1][3][12]  (.D(\input_filter[1][3] [12]), .CK(n_58_15), 
      .Q(\buffer[15][1][3] [12]), .QN());
   DFF_X1 \buffer_reg[15][1][3][11]  (.D(\input_filter[1][3] [11]), .CK(n_58_15), 
      .Q(\buffer[15][1][3] [11]), .QN());
   DFF_X1 \buffer_reg[15][1][3][10]  (.D(\input_filter[1][3] [10]), .CK(n_58_15), 
      .Q(\buffer[15][1][3] [10]), .QN());
   DFF_X1 \buffer_reg[15][1][3][9]  (.D(\input_filter[1][3] [9]), .CK(n_58_15), 
      .Q(\buffer[15][1][3] [9]), .QN());
   DFF_X1 \buffer_reg[15][1][3][8]  (.D(\input_filter[1][3] [8]), .CK(n_58_15), 
      .Q(\buffer[15][1][3] [8]), .QN());
   DFF_X1 \buffer_reg[15][1][3][7]  (.D(\input_filter[1][3] [7]), .CK(n_58_15), 
      .Q(\buffer[15][1][3] [7]), .QN());
   DFF_X1 \buffer_reg[15][1][3][6]  (.D(\input_filter[1][3] [6]), .CK(n_58_15), 
      .Q(\buffer[15][1][3] [6]), .QN());
   DFF_X1 \buffer_reg[15][1][3][5]  (.D(\input_filter[1][3] [5]), .CK(n_58_15), 
      .Q(\buffer[15][1][3] [5]), .QN());
   DFF_X1 \buffer_reg[15][1][3][4]  (.D(\input_filter[1][3] [4]), .CK(n_58_15), 
      .Q(\buffer[15][1][3] [4]), .QN());
   DFF_X1 \buffer_reg[15][1][3][3]  (.D(\input_filter[1][3] [3]), .CK(n_58_15), 
      .Q(\buffer[15][1][3] [3]), .QN());
   DFF_X1 \buffer_reg[15][1][3][2]  (.D(\input_filter[1][3] [2]), .CK(n_58_15), 
      .Q(\buffer[15][1][3] [2]), .QN());
   DFF_X1 \buffer_reg[15][1][3][1]  (.D(\input_filter[1][3] [1]), .CK(n_58_15), 
      .Q(\buffer[15][1][3] [1]), .QN());
   DFF_X1 \buffer_reg[15][1][3][0]  (.D(\input_filter[1][3] [0]), .CK(n_58_15), 
      .Q(\buffer[15][1][3] [0]), .QN());
   DFF_X1 \buffer_reg[5][0][2][15]  (.D(\input_filter[0][2] [15]), .CK(n_58_5), 
      .Q(\buffer[5][0][2] [15]), .QN());
   DFF_X1 \buffer_reg[5][0][2][14]  (.D(\input_filter[0][2] [14]), .CK(n_58_5), 
      .Q(\buffer[5][0][2] [14]), .QN());
   DFF_X1 \buffer_reg[5][0][2][13]  (.D(\input_filter[0][2] [13]), .CK(n_58_5), 
      .Q(\buffer[5][0][2] [13]), .QN());
   DFF_X1 \buffer_reg[5][0][2][12]  (.D(\input_filter[0][2] [12]), .CK(n_58_5), 
      .Q(\buffer[5][0][2] [12]), .QN());
   DFF_X1 \buffer_reg[5][0][2][11]  (.D(\input_filter[0][2] [11]), .CK(n_58_5), 
      .Q(\buffer[5][0][2] [11]), .QN());
   DFF_X1 \buffer_reg[5][0][2][10]  (.D(\input_filter[0][2] [10]), .CK(n_58_5), 
      .Q(\buffer[5][0][2] [10]), .QN());
   DFF_X1 \buffer_reg[5][0][2][9]  (.D(\input_filter[0][2] [9]), .CK(n_58_5), 
      .Q(\buffer[5][0][2] [9]), .QN());
   DFF_X1 \buffer_reg[5][0][2][8]  (.D(\input_filter[0][2] [8]), .CK(n_58_5), 
      .Q(\buffer[5][0][2] [8]), .QN());
   DFF_X1 \buffer_reg[5][0][2][7]  (.D(\input_filter[0][2] [7]), .CK(n_58_5), 
      .Q(\buffer[5][0][2] [7]), .QN());
   DFF_X1 \buffer_reg[5][0][2][6]  (.D(\input_filter[0][2] [6]), .CK(n_58_5), 
      .Q(\buffer[5][0][2] [6]), .QN());
   DFF_X1 \buffer_reg[5][0][2][5]  (.D(\input_filter[0][2] [5]), .CK(n_58_5), 
      .Q(\buffer[5][0][2] [5]), .QN());
   DFF_X1 \buffer_reg[5][0][2][4]  (.D(\input_filter[0][2] [4]), .CK(n_58_5), 
      .Q(\buffer[5][0][2] [4]), .QN());
   DFF_X1 \buffer_reg[5][0][2][3]  (.D(\input_filter[0][2] [3]), .CK(n_58_5), 
      .Q(\buffer[5][0][2] [3]), .QN());
   DFF_X1 \buffer_reg[5][0][2][2]  (.D(\input_filter[0][2] [2]), .CK(n_58_5), 
      .Q(\buffer[5][0][2] [2]), .QN());
   DFF_X1 \buffer_reg[5][0][2][1]  (.D(\input_filter[0][2] [1]), .CK(n_58_5), 
      .Q(\buffer[5][0][2] [1]), .QN());
   DFF_X1 \buffer_reg[5][0][2][0]  (.D(\input_filter[0][2] [0]), .CK(n_58_5), 
      .Q(\buffer[5][0][2] [0]), .QN());
   DFF_X1 \buffer_reg[4][0][2][15]  (.D(\input_filter[0][2] [15]), .CK(n_58_4), 
      .Q(\buffer[4][0][2] [15]), .QN());
   DFF_X1 \buffer_reg[4][0][2][14]  (.D(\input_filter[0][2] [14]), .CK(n_58_4), 
      .Q(\buffer[4][0][2] [14]), .QN());
   DFF_X1 \buffer_reg[4][0][2][13]  (.D(\input_filter[0][2] [13]), .CK(n_58_4), 
      .Q(\buffer[4][0][2] [13]), .QN());
   DFF_X1 \buffer_reg[4][0][2][12]  (.D(\input_filter[0][2] [12]), .CK(n_58_4), 
      .Q(\buffer[4][0][2] [12]), .QN());
   DFF_X1 \buffer_reg[4][0][2][11]  (.D(\input_filter[0][2] [11]), .CK(n_58_4), 
      .Q(\buffer[4][0][2] [11]), .QN());
   DFF_X1 \buffer_reg[4][0][2][10]  (.D(\input_filter[0][2] [10]), .CK(n_58_4), 
      .Q(\buffer[4][0][2] [10]), .QN());
   DFF_X1 \buffer_reg[4][0][2][9]  (.D(\input_filter[0][2] [9]), .CK(n_58_4), 
      .Q(\buffer[4][0][2] [9]), .QN());
   DFF_X1 \buffer_reg[4][0][2][8]  (.D(\input_filter[0][2] [8]), .CK(n_58_4), 
      .Q(\buffer[4][0][2] [8]), .QN());
   DFF_X1 \buffer_reg[4][0][2][7]  (.D(\input_filter[0][2] [7]), .CK(n_58_4), 
      .Q(\buffer[4][0][2] [7]), .QN());
   DFF_X1 \buffer_reg[4][0][2][6]  (.D(\input_filter[0][2] [6]), .CK(n_58_4), 
      .Q(\buffer[4][0][2] [6]), .QN());
   DFF_X1 \buffer_reg[4][0][2][5]  (.D(\input_filter[0][2] [5]), .CK(n_58_4), 
      .Q(\buffer[4][0][2] [5]), .QN());
   DFF_X1 \buffer_reg[4][0][2][4]  (.D(\input_filter[0][2] [4]), .CK(n_58_4), 
      .Q(\buffer[4][0][2] [4]), .QN());
   DFF_X1 \buffer_reg[4][0][2][3]  (.D(\input_filter[0][2] [3]), .CK(n_58_4), 
      .Q(\buffer[4][0][2] [3]), .QN());
   DFF_X1 \buffer_reg[4][0][2][2]  (.D(\input_filter[0][2] [2]), .CK(n_58_4), 
      .Q(\buffer[4][0][2] [2]), .QN());
   DFF_X1 \buffer_reg[4][0][2][1]  (.D(\input_filter[0][2] [1]), .CK(n_58_4), 
      .Q(\buffer[4][0][2] [1]), .QN());
   DFF_X1 \buffer_reg[4][0][2][0]  (.D(\input_filter[0][2] [0]), .CK(n_58_4), 
      .Q(\buffer[4][0][2] [0]), .QN());
   DFF_X1 \buffer_reg[3][0][2][15]  (.D(\input_filter[0][2] [15]), .CK(n_58_3), 
      .Q(\buffer[3][0][2] [15]), .QN());
   DFF_X1 \buffer_reg[3][0][2][14]  (.D(\input_filter[0][2] [14]), .CK(n_58_3), 
      .Q(\buffer[3][0][2] [14]), .QN());
   DFF_X1 \buffer_reg[3][0][2][13]  (.D(\input_filter[0][2] [13]), .CK(n_58_3), 
      .Q(\buffer[3][0][2] [13]), .QN());
   DFF_X1 \buffer_reg[3][0][2][12]  (.D(\input_filter[0][2] [12]), .CK(n_58_3), 
      .Q(\buffer[3][0][2] [12]), .QN());
   DFF_X1 \buffer_reg[3][0][2][11]  (.D(\input_filter[0][2] [11]), .CK(n_58_3), 
      .Q(\buffer[3][0][2] [11]), .QN());
   DFF_X1 \buffer_reg[3][0][2][10]  (.D(\input_filter[0][2] [10]), .CK(n_58_3), 
      .Q(\buffer[3][0][2] [10]), .QN());
   DFF_X1 \buffer_reg[3][0][2][9]  (.D(\input_filter[0][2] [9]), .CK(n_58_3), 
      .Q(\buffer[3][0][2] [9]), .QN());
   DFF_X1 \buffer_reg[3][0][2][8]  (.D(\input_filter[0][2] [8]), .CK(n_58_3), 
      .Q(\buffer[3][0][2] [8]), .QN());
   DFF_X1 \buffer_reg[3][0][2][7]  (.D(\input_filter[0][2] [7]), .CK(n_58_3), 
      .Q(\buffer[3][0][2] [7]), .QN());
   DFF_X1 \buffer_reg[3][0][2][6]  (.D(\input_filter[0][2] [6]), .CK(n_58_3), 
      .Q(\buffer[3][0][2] [6]), .QN());
   DFF_X1 \buffer_reg[3][0][2][5]  (.D(\input_filter[0][2] [5]), .CK(n_58_3), 
      .Q(\buffer[3][0][2] [5]), .QN());
   DFF_X1 \buffer_reg[3][0][2][4]  (.D(\input_filter[0][2] [4]), .CK(n_58_3), 
      .Q(\buffer[3][0][2] [4]), .QN());
   DFF_X1 \buffer_reg[3][0][2][3]  (.D(\input_filter[0][2] [3]), .CK(n_58_3), 
      .Q(\buffer[3][0][2] [3]), .QN());
   DFF_X1 \buffer_reg[3][0][2][2]  (.D(\input_filter[0][2] [2]), .CK(n_58_3), 
      .Q(\buffer[3][0][2] [2]), .QN());
   DFF_X1 \buffer_reg[3][0][2][1]  (.D(\input_filter[0][2] [1]), .CK(n_58_3), 
      .Q(\buffer[3][0][2] [1]), .QN());
   DFF_X1 \buffer_reg[3][0][2][0]  (.D(\input_filter[0][2] [0]), .CK(n_58_3), 
      .Q(\buffer[3][0][2] [0]), .QN());
   DFF_X1 \buffer_reg[2][0][2][15]  (.D(\input_filter[0][2] [15]), .CK(n_58_2), 
      .Q(\buffer[2][0][2] [15]), .QN());
   DFF_X1 \buffer_reg[2][0][2][14]  (.D(\input_filter[0][2] [14]), .CK(n_58_2), 
      .Q(\buffer[2][0][2] [14]), .QN());
   DFF_X1 \buffer_reg[2][0][2][13]  (.D(\input_filter[0][2] [13]), .CK(n_58_2), 
      .Q(\buffer[2][0][2] [13]), .QN());
   DFF_X1 \buffer_reg[2][0][2][12]  (.D(\input_filter[0][2] [12]), .CK(n_58_2), 
      .Q(\buffer[2][0][2] [12]), .QN());
   DFF_X1 \buffer_reg[2][0][2][11]  (.D(\input_filter[0][2] [11]), .CK(n_58_2), 
      .Q(\buffer[2][0][2] [11]), .QN());
   DFF_X1 \buffer_reg[2][0][2][10]  (.D(\input_filter[0][2] [10]), .CK(n_58_2), 
      .Q(\buffer[2][0][2] [10]), .QN());
   DFF_X1 \buffer_reg[2][0][2][9]  (.D(\input_filter[0][2] [9]), .CK(n_58_2), 
      .Q(\buffer[2][0][2] [9]), .QN());
   DFF_X1 \buffer_reg[2][0][2][8]  (.D(\input_filter[0][2] [8]), .CK(n_58_2), 
      .Q(\buffer[2][0][2] [8]), .QN());
   DFF_X1 \buffer_reg[2][0][2][7]  (.D(\input_filter[0][2] [7]), .CK(n_58_2), 
      .Q(\buffer[2][0][2] [7]), .QN());
   DFF_X1 \buffer_reg[2][0][2][6]  (.D(\input_filter[0][2] [6]), .CK(n_58_2), 
      .Q(\buffer[2][0][2] [6]), .QN());
   DFF_X1 \buffer_reg[2][0][2][5]  (.D(\input_filter[0][2] [5]), .CK(n_58_2), 
      .Q(\buffer[2][0][2] [5]), .QN());
   DFF_X1 \buffer_reg[2][0][2][4]  (.D(\input_filter[0][2] [4]), .CK(n_58_2), 
      .Q(\buffer[2][0][2] [4]), .QN());
   DFF_X1 \buffer_reg[2][0][2][3]  (.D(\input_filter[0][2] [3]), .CK(n_58_2), 
      .Q(\buffer[2][0][2] [3]), .QN());
   DFF_X1 \buffer_reg[2][0][2][2]  (.D(\input_filter[0][2] [2]), .CK(n_58_2), 
      .Q(\buffer[2][0][2] [2]), .QN());
   DFF_X1 \buffer_reg[2][0][2][1]  (.D(\input_filter[0][2] [1]), .CK(n_58_2), 
      .Q(\buffer[2][0][2] [1]), .QN());
   DFF_X1 \buffer_reg[2][0][2][0]  (.D(\input_filter[0][2] [0]), .CK(n_58_2), 
      .Q(\buffer[2][0][2] [0]), .QN());
   DFF_X1 \buffer_reg[0][0][3][15]  (.D(\input_filter[0][3] [15]), .CK(n_58_0), 
      .Q(\buffer[0][0][3] [15]), .QN());
   DFF_X1 \buffer_reg[0][0][3][14]  (.D(\input_filter[0][3] [14]), .CK(n_58_0), 
      .Q(\buffer[0][0][3] [14]), .QN());
   DFF_X1 \buffer_reg[0][0][3][13]  (.D(\input_filter[0][3] [13]), .CK(n_58_0), 
      .Q(\buffer[0][0][3] [13]), .QN());
   DFF_X1 \buffer_reg[0][0][3][12]  (.D(\input_filter[0][3] [12]), .CK(n_58_0), 
      .Q(\buffer[0][0][3] [12]), .QN());
   DFF_X1 \buffer_reg[0][0][3][11]  (.D(\input_filter[0][3] [11]), .CK(n_58_0), 
      .Q(\buffer[0][0][3] [11]), .QN());
   DFF_X1 \buffer_reg[0][0][3][10]  (.D(\input_filter[0][3] [10]), .CK(n_58_0), 
      .Q(\buffer[0][0][3] [10]), .QN());
   DFF_X1 \buffer_reg[0][0][3][9]  (.D(\input_filter[0][3] [9]), .CK(n_58_0), 
      .Q(\buffer[0][0][3] [9]), .QN());
   DFF_X1 \buffer_reg[0][0][3][8]  (.D(\input_filter[0][3] [8]), .CK(n_58_0), 
      .Q(\buffer[0][0][3] [8]), .QN());
   DFF_X1 \buffer_reg[0][0][3][7]  (.D(\input_filter[0][3] [7]), .CK(n_58_0), 
      .Q(\buffer[0][0][3] [7]), .QN());
   DFF_X1 \buffer_reg[0][0][3][6]  (.D(\input_filter[0][3] [6]), .CK(n_58_0), 
      .Q(\buffer[0][0][3] [6]), .QN());
   DFF_X1 \buffer_reg[0][0][3][5]  (.D(\input_filter[0][3] [5]), .CK(n_58_0), 
      .Q(\buffer[0][0][3] [5]), .QN());
   DFF_X1 \buffer_reg[0][0][3][4]  (.D(\input_filter[0][3] [4]), .CK(n_58_0), 
      .Q(\buffer[0][0][3] [4]), .QN());
   DFF_X1 \buffer_reg[0][0][3][3]  (.D(\input_filter[0][3] [3]), .CK(n_58_0), 
      .Q(\buffer[0][0][3] [3]), .QN());
   DFF_X1 \buffer_reg[0][0][3][2]  (.D(\input_filter[0][3] [2]), .CK(n_58_0), 
      .Q(\buffer[0][0][3] [2]), .QN());
   DFF_X1 \buffer_reg[0][0][3][1]  (.D(\input_filter[0][3] [1]), .CK(n_58_0), 
      .Q(\buffer[0][0][3] [1]), .QN());
   DFF_X1 \buffer_reg[0][0][3][0]  (.D(\input_filter[0][3] [0]), .CK(n_58_0), 
      .Q(\buffer[0][0][3] [0]), .QN());
   DFF_X1 \buffer_reg[1][0][2][15]  (.D(\input_filter[0][2] [15]), .CK(n_58_1), 
      .Q(\buffer[1][0][2] [15]), .QN());
   DFF_X1 \buffer_reg[1][0][2][14]  (.D(\input_filter[0][2] [14]), .CK(n_58_1), 
      .Q(\buffer[1][0][2] [14]), .QN());
   DFF_X1 \buffer_reg[1][0][2][13]  (.D(\input_filter[0][2] [13]), .CK(n_58_1), 
      .Q(\buffer[1][0][2] [13]), .QN());
   DFF_X1 \buffer_reg[1][0][2][12]  (.D(\input_filter[0][2] [12]), .CK(n_58_1), 
      .Q(\buffer[1][0][2] [12]), .QN());
   DFF_X1 \buffer_reg[1][0][2][11]  (.D(\input_filter[0][2] [11]), .CK(n_58_1), 
      .Q(\buffer[1][0][2] [11]), .QN());
   DFF_X1 \buffer_reg[1][0][2][10]  (.D(\input_filter[0][2] [10]), .CK(n_58_1), 
      .Q(\buffer[1][0][2] [10]), .QN());
   DFF_X1 \buffer_reg[1][0][2][9]  (.D(\input_filter[0][2] [9]), .CK(n_58_1), 
      .Q(\buffer[1][0][2] [9]), .QN());
   DFF_X1 \buffer_reg[1][0][2][8]  (.D(\input_filter[0][2] [8]), .CK(n_58_1), 
      .Q(\buffer[1][0][2] [8]), .QN());
   DFF_X1 \buffer_reg[1][0][2][7]  (.D(\input_filter[0][2] [7]), .CK(n_58_1), 
      .Q(\buffer[1][0][2] [7]), .QN());
   DFF_X1 \buffer_reg[1][0][2][6]  (.D(\input_filter[0][2] [6]), .CK(n_58_1), 
      .Q(\buffer[1][0][2] [6]), .QN());
   DFF_X1 \buffer_reg[1][0][2][5]  (.D(\input_filter[0][2] [5]), .CK(n_58_1), 
      .Q(\buffer[1][0][2] [5]), .QN());
   DFF_X1 \buffer_reg[1][0][2][4]  (.D(\input_filter[0][2] [4]), .CK(n_58_1), 
      .Q(\buffer[1][0][2] [4]), .QN());
   DFF_X1 \buffer_reg[1][0][2][3]  (.D(\input_filter[0][2] [3]), .CK(n_58_1), 
      .Q(\buffer[1][0][2] [3]), .QN());
   DFF_X1 \buffer_reg[1][0][2][2]  (.D(\input_filter[0][2] [2]), .CK(n_58_1), 
      .Q(\buffer[1][0][2] [2]), .QN());
   DFF_X1 \buffer_reg[1][0][2][1]  (.D(\input_filter[0][2] [1]), .CK(n_58_1), 
      .Q(\buffer[1][0][2] [1]), .QN());
   DFF_X1 \buffer_reg[1][0][2][0]  (.D(\input_filter[0][2] [0]), .CK(n_58_1), 
      .Q(\buffer[1][0][2] [0]), .QN());
   DFF_X1 \buffer_reg[14][0][2][15]  (.D(\input_filter[0][2] [15]), .CK(n_58_14), 
      .Q(\buffer[14][0][2] [15]), .QN());
   DFF_X1 \buffer_reg[14][0][2][14]  (.D(\input_filter[0][2] [14]), .CK(n_58_14), 
      .Q(\buffer[14][0][2] [14]), .QN());
   DFF_X1 \buffer_reg[14][0][2][13]  (.D(\input_filter[0][2] [13]), .CK(n_58_14), 
      .Q(\buffer[14][0][2] [13]), .QN());
   DFF_X1 \buffer_reg[14][0][2][12]  (.D(\input_filter[0][2] [12]), .CK(n_58_14), 
      .Q(\buffer[14][0][2] [12]), .QN());
   DFF_X1 \buffer_reg[14][0][2][11]  (.D(\input_filter[0][2] [11]), .CK(n_58_14), 
      .Q(\buffer[14][0][2] [11]), .QN());
   DFF_X1 \buffer_reg[14][0][2][10]  (.D(\input_filter[0][2] [10]), .CK(n_58_14), 
      .Q(\buffer[14][0][2] [10]), .QN());
   DFF_X1 \buffer_reg[14][0][2][9]  (.D(\input_filter[0][2] [9]), .CK(n_58_14), 
      .Q(\buffer[14][0][2] [9]), .QN());
   DFF_X1 \buffer_reg[14][0][2][8]  (.D(\input_filter[0][2] [8]), .CK(n_58_14), 
      .Q(\buffer[14][0][2] [8]), .QN());
   DFF_X1 \buffer_reg[14][0][2][7]  (.D(\input_filter[0][2] [7]), .CK(n_58_14), 
      .Q(\buffer[14][0][2] [7]), .QN());
   DFF_X1 \buffer_reg[14][0][2][6]  (.D(\input_filter[0][2] [6]), .CK(n_58_14), 
      .Q(\buffer[14][0][2] [6]), .QN());
   DFF_X1 \buffer_reg[14][0][2][5]  (.D(\input_filter[0][2] [5]), .CK(n_58_14), 
      .Q(\buffer[14][0][2] [5]), .QN());
   DFF_X1 \buffer_reg[14][0][2][4]  (.D(\input_filter[0][2] [4]), .CK(n_58_14), 
      .Q(\buffer[14][0][2] [4]), .QN());
   DFF_X1 \buffer_reg[14][0][2][3]  (.D(\input_filter[0][2] [3]), .CK(n_58_14), 
      .Q(\buffer[14][0][2] [3]), .QN());
   DFF_X1 \buffer_reg[14][0][2][2]  (.D(\input_filter[0][2] [2]), .CK(n_58_14), 
      .Q(\buffer[14][0][2] [2]), .QN());
   DFF_X1 \buffer_reg[14][0][2][1]  (.D(\input_filter[0][2] [1]), .CK(n_58_14), 
      .Q(\buffer[14][0][2] [1]), .QN());
   DFF_X1 \buffer_reg[14][0][2][0]  (.D(\input_filter[0][2] [0]), .CK(n_58_14), 
      .Q(\buffer[14][0][2] [0]), .QN());
   DFF_X1 \buffer_reg[13][0][2][15]  (.D(\input_filter[0][2] [15]), .CK(n_58_13), 
      .Q(\buffer[13][0][2] [15]), .QN());
   DFF_X1 \buffer_reg[13][0][2][14]  (.D(\input_filter[0][2] [14]), .CK(n_58_13), 
      .Q(\buffer[13][0][2] [14]), .QN());
   DFF_X1 \buffer_reg[13][0][2][13]  (.D(\input_filter[0][2] [13]), .CK(n_58_13), 
      .Q(\buffer[13][0][2] [13]), .QN());
   DFF_X1 \buffer_reg[13][0][2][12]  (.D(\input_filter[0][2] [12]), .CK(n_58_13), 
      .Q(\buffer[13][0][2] [12]), .QN());
   DFF_X1 \buffer_reg[13][0][2][11]  (.D(\input_filter[0][2] [11]), .CK(n_58_13), 
      .Q(\buffer[13][0][2] [11]), .QN());
   DFF_X1 \buffer_reg[13][0][2][10]  (.D(\input_filter[0][2] [10]), .CK(n_58_13), 
      .Q(\buffer[13][0][2] [10]), .QN());
   DFF_X1 \buffer_reg[13][0][2][9]  (.D(\input_filter[0][2] [9]), .CK(n_58_13), 
      .Q(\buffer[13][0][2] [9]), .QN());
   DFF_X1 \buffer_reg[13][0][2][8]  (.D(\input_filter[0][2] [8]), .CK(n_58_13), 
      .Q(\buffer[13][0][2] [8]), .QN());
   DFF_X1 \buffer_reg[13][0][2][7]  (.D(\input_filter[0][2] [7]), .CK(n_58_13), 
      .Q(\buffer[13][0][2] [7]), .QN());
   DFF_X1 \buffer_reg[13][0][2][6]  (.D(\input_filter[0][2] [6]), .CK(n_58_13), 
      .Q(\buffer[13][0][2] [6]), .QN());
   DFF_X1 \buffer_reg[13][0][2][5]  (.D(\input_filter[0][2] [5]), .CK(n_58_13), 
      .Q(\buffer[13][0][2] [5]), .QN());
   DFF_X1 \buffer_reg[13][0][2][4]  (.D(\input_filter[0][2] [4]), .CK(n_58_13), 
      .Q(\buffer[13][0][2] [4]), .QN());
   DFF_X1 \buffer_reg[13][0][2][3]  (.D(\input_filter[0][2] [3]), .CK(n_58_13), 
      .Q(\buffer[13][0][2] [3]), .QN());
   DFF_X1 \buffer_reg[13][0][2][2]  (.D(\input_filter[0][2] [2]), .CK(n_58_13), 
      .Q(\buffer[13][0][2] [2]), .QN());
   DFF_X1 \buffer_reg[13][0][2][1]  (.D(\input_filter[0][2] [1]), .CK(n_58_13), 
      .Q(\buffer[13][0][2] [1]), .QN());
   DFF_X1 \buffer_reg[13][0][2][0]  (.D(\input_filter[0][2] [0]), .CK(n_58_13), 
      .Q(\buffer[13][0][2] [0]), .QN());
   DFF_X1 \buffer_reg[12][0][2][15]  (.D(\input_filter[0][2] [15]), .CK(n_58_12), 
      .Q(\buffer[12][0][2] [15]), .QN());
   DFF_X1 \buffer_reg[12][0][2][14]  (.D(\input_filter[0][2] [14]), .CK(n_58_12), 
      .Q(\buffer[12][0][2] [14]), .QN());
   DFF_X1 \buffer_reg[12][0][2][13]  (.D(\input_filter[0][2] [13]), .CK(n_58_12), 
      .Q(\buffer[12][0][2] [13]), .QN());
   DFF_X1 \buffer_reg[12][0][2][12]  (.D(\input_filter[0][2] [12]), .CK(n_58_12), 
      .Q(\buffer[12][0][2] [12]), .QN());
   DFF_X1 \buffer_reg[12][0][2][11]  (.D(\input_filter[0][2] [11]), .CK(n_58_12), 
      .Q(\buffer[12][0][2] [11]), .QN());
   DFF_X1 \buffer_reg[12][0][2][10]  (.D(\input_filter[0][2] [10]), .CK(n_58_12), 
      .Q(\buffer[12][0][2] [10]), .QN());
   DFF_X1 \buffer_reg[12][0][2][9]  (.D(\input_filter[0][2] [9]), .CK(n_58_12), 
      .Q(\buffer[12][0][2] [9]), .QN());
   DFF_X1 \buffer_reg[12][0][2][8]  (.D(\input_filter[0][2] [8]), .CK(n_58_12), 
      .Q(\buffer[12][0][2] [8]), .QN());
   DFF_X1 \buffer_reg[12][0][2][7]  (.D(\input_filter[0][2] [7]), .CK(n_58_12), 
      .Q(\buffer[12][0][2] [7]), .QN());
   DFF_X1 \buffer_reg[12][0][2][6]  (.D(\input_filter[0][2] [6]), .CK(n_58_12), 
      .Q(\buffer[12][0][2] [6]), .QN());
   DFF_X1 \buffer_reg[12][0][2][5]  (.D(\input_filter[0][2] [5]), .CK(n_58_12), 
      .Q(\buffer[12][0][2] [5]), .QN());
   DFF_X1 \buffer_reg[12][0][2][4]  (.D(\input_filter[0][2] [4]), .CK(n_58_12), 
      .Q(\buffer[12][0][2] [4]), .QN());
   DFF_X1 \buffer_reg[12][0][2][3]  (.D(\input_filter[0][2] [3]), .CK(n_58_12), 
      .Q(\buffer[12][0][2] [3]), .QN());
   DFF_X1 \buffer_reg[12][0][2][2]  (.D(\input_filter[0][2] [2]), .CK(n_58_12), 
      .Q(\buffer[12][0][2] [2]), .QN());
   DFF_X1 \buffer_reg[12][0][2][1]  (.D(\input_filter[0][2] [1]), .CK(n_58_12), 
      .Q(\buffer[12][0][2] [1]), .QN());
   DFF_X1 \buffer_reg[12][0][2][0]  (.D(\input_filter[0][2] [0]), .CK(n_58_12), 
      .Q(\buffer[12][0][2] [0]), .QN());
   DFF_X1 \buffer_reg[11][0][2][15]  (.D(\input_filter[0][2] [15]), .CK(n_58_11), 
      .Q(\buffer[11][0][2] [15]), .QN());
   DFF_X1 \buffer_reg[11][0][2][14]  (.D(\input_filter[0][2] [14]), .CK(n_58_11), 
      .Q(\buffer[11][0][2] [14]), .QN());
   DFF_X1 \buffer_reg[11][0][2][13]  (.D(\input_filter[0][2] [13]), .CK(n_58_11), 
      .Q(\buffer[11][0][2] [13]), .QN());
   DFF_X1 \buffer_reg[11][0][2][12]  (.D(\input_filter[0][2] [12]), .CK(n_58_11), 
      .Q(\buffer[11][0][2] [12]), .QN());
   DFF_X1 \buffer_reg[11][0][2][11]  (.D(\input_filter[0][2] [11]), .CK(n_58_11), 
      .Q(\buffer[11][0][2] [11]), .QN());
   DFF_X1 \buffer_reg[11][0][2][10]  (.D(\input_filter[0][2] [10]), .CK(n_58_11), 
      .Q(\buffer[11][0][2] [10]), .QN());
   DFF_X1 \buffer_reg[11][0][2][9]  (.D(\input_filter[0][2] [9]), .CK(n_58_11), 
      .Q(\buffer[11][0][2] [9]), .QN());
   DFF_X1 \buffer_reg[11][0][2][8]  (.D(\input_filter[0][2] [8]), .CK(n_58_11), 
      .Q(\buffer[11][0][2] [8]), .QN());
   DFF_X1 \buffer_reg[11][0][2][7]  (.D(\input_filter[0][2] [7]), .CK(n_58_11), 
      .Q(\buffer[11][0][2] [7]), .QN());
   DFF_X1 \buffer_reg[11][0][2][6]  (.D(\input_filter[0][2] [6]), .CK(n_58_11), 
      .Q(\buffer[11][0][2] [6]), .QN());
   DFF_X1 \buffer_reg[11][0][2][5]  (.D(\input_filter[0][2] [5]), .CK(n_58_11), 
      .Q(\buffer[11][0][2] [5]), .QN());
   DFF_X1 \buffer_reg[11][0][2][4]  (.D(\input_filter[0][2] [4]), .CK(n_58_11), 
      .Q(\buffer[11][0][2] [4]), .QN());
   DFF_X1 \buffer_reg[11][0][2][3]  (.D(\input_filter[0][2] [3]), .CK(n_58_11), 
      .Q(\buffer[11][0][2] [3]), .QN());
   DFF_X1 \buffer_reg[11][0][2][2]  (.D(\input_filter[0][2] [2]), .CK(n_58_11), 
      .Q(\buffer[11][0][2] [2]), .QN());
   DFF_X1 \buffer_reg[11][0][2][1]  (.D(\input_filter[0][2] [1]), .CK(n_58_11), 
      .Q(\buffer[11][0][2] [1]), .QN());
   DFF_X1 \buffer_reg[11][0][2][0]  (.D(\input_filter[0][2] [0]), .CK(n_58_11), 
      .Q(\buffer[11][0][2] [0]), .QN());
   DFF_X1 \buffer_reg[10][0][2][15]  (.D(\input_filter[0][2] [15]), .CK(n_58_10), 
      .Q(\buffer[10][0][2] [15]), .QN());
   DFF_X1 \buffer_reg[10][0][2][14]  (.D(\input_filter[0][2] [14]), .CK(n_58_10), 
      .Q(\buffer[10][0][2] [14]), .QN());
   DFF_X1 \buffer_reg[10][0][2][13]  (.D(\input_filter[0][2] [13]), .CK(n_58_10), 
      .Q(\buffer[10][0][2] [13]), .QN());
   DFF_X1 \buffer_reg[10][0][2][12]  (.D(\input_filter[0][2] [12]), .CK(n_58_10), 
      .Q(\buffer[10][0][2] [12]), .QN());
   DFF_X1 \buffer_reg[10][0][2][11]  (.D(\input_filter[0][2] [11]), .CK(n_58_10), 
      .Q(\buffer[10][0][2] [11]), .QN());
   DFF_X1 \buffer_reg[10][0][2][10]  (.D(\input_filter[0][2] [10]), .CK(n_58_10), 
      .Q(\buffer[10][0][2] [10]), .QN());
   DFF_X1 \buffer_reg[10][0][2][9]  (.D(\input_filter[0][2] [9]), .CK(n_58_10), 
      .Q(\buffer[10][0][2] [9]), .QN());
   DFF_X1 \buffer_reg[10][0][2][8]  (.D(\input_filter[0][2] [8]), .CK(n_58_10), 
      .Q(\buffer[10][0][2] [8]), .QN());
   DFF_X1 \buffer_reg[10][0][2][7]  (.D(\input_filter[0][2] [7]), .CK(n_58_10), 
      .Q(\buffer[10][0][2] [7]), .QN());
   DFF_X1 \buffer_reg[10][0][2][6]  (.D(\input_filter[0][2] [6]), .CK(n_58_10), 
      .Q(\buffer[10][0][2] [6]), .QN());
   DFF_X1 \buffer_reg[10][0][2][5]  (.D(\input_filter[0][2] [5]), .CK(n_58_10), 
      .Q(\buffer[10][0][2] [5]), .QN());
   DFF_X1 \buffer_reg[10][0][2][4]  (.D(\input_filter[0][2] [4]), .CK(n_58_10), 
      .Q(\buffer[10][0][2] [4]), .QN());
   DFF_X1 \buffer_reg[10][0][2][3]  (.D(\input_filter[0][2] [3]), .CK(n_58_10), 
      .Q(\buffer[10][0][2] [3]), .QN());
   DFF_X1 \buffer_reg[10][0][2][2]  (.D(\input_filter[0][2] [2]), .CK(n_58_10), 
      .Q(\buffer[10][0][2] [2]), .QN());
   DFF_X1 \buffer_reg[10][0][2][1]  (.D(\input_filter[0][2] [1]), .CK(n_58_10), 
      .Q(\buffer[10][0][2] [1]), .QN());
   DFF_X1 \buffer_reg[10][0][2][0]  (.D(\input_filter[0][2] [0]), .CK(n_58_10), 
      .Q(\buffer[10][0][2] [0]), .QN());
   DFF_X1 \buffer_reg[9][0][2][15]  (.D(\input_filter[0][2] [15]), .CK(n_58_9), 
      .Q(\buffer[9][0][2] [15]), .QN());
   DFF_X1 \buffer_reg[9][0][2][14]  (.D(\input_filter[0][2] [14]), .CK(n_58_9), 
      .Q(\buffer[9][0][2] [14]), .QN());
   DFF_X1 \buffer_reg[9][0][2][13]  (.D(\input_filter[0][2] [13]), .CK(n_58_9), 
      .Q(\buffer[9][0][2] [13]), .QN());
   DFF_X1 \buffer_reg[9][0][2][12]  (.D(\input_filter[0][2] [12]), .CK(n_58_9), 
      .Q(\buffer[9][0][2] [12]), .QN());
   DFF_X1 \buffer_reg[9][0][2][11]  (.D(\input_filter[0][2] [11]), .CK(n_58_9), 
      .Q(\buffer[9][0][2] [11]), .QN());
   DFF_X1 \buffer_reg[9][0][2][10]  (.D(\input_filter[0][2] [10]), .CK(n_58_9), 
      .Q(\buffer[9][0][2] [10]), .QN());
   DFF_X1 \buffer_reg[9][0][2][9]  (.D(\input_filter[0][2] [9]), .CK(n_58_9), 
      .Q(\buffer[9][0][2] [9]), .QN());
   DFF_X1 \buffer_reg[9][0][2][8]  (.D(\input_filter[0][2] [8]), .CK(n_58_9), 
      .Q(\buffer[9][0][2] [8]), .QN());
   DFF_X1 \buffer_reg[9][0][2][7]  (.D(\input_filter[0][2] [7]), .CK(n_58_9), 
      .Q(\buffer[9][0][2] [7]), .QN());
   DFF_X1 \buffer_reg[9][0][2][6]  (.D(\input_filter[0][2] [6]), .CK(n_58_9), 
      .Q(\buffer[9][0][2] [6]), .QN());
   DFF_X1 \buffer_reg[9][0][2][5]  (.D(\input_filter[0][2] [5]), .CK(n_58_9), 
      .Q(\buffer[9][0][2] [5]), .QN());
   DFF_X1 \buffer_reg[9][0][2][4]  (.D(\input_filter[0][2] [4]), .CK(n_58_9), 
      .Q(\buffer[9][0][2] [4]), .QN());
   DFF_X1 \buffer_reg[9][0][2][3]  (.D(\input_filter[0][2] [3]), .CK(n_58_9), 
      .Q(\buffer[9][0][2] [3]), .QN());
   DFF_X1 \buffer_reg[9][0][2][2]  (.D(\input_filter[0][2] [2]), .CK(n_58_9), 
      .Q(\buffer[9][0][2] [2]), .QN());
   DFF_X1 \buffer_reg[9][0][2][1]  (.D(\input_filter[0][2] [1]), .CK(n_58_9), 
      .Q(\buffer[9][0][2] [1]), .QN());
   DFF_X1 \buffer_reg[9][0][2][0]  (.D(\input_filter[0][2] [0]), .CK(n_58_9), 
      .Q(\buffer[9][0][2] [0]), .QN());
   DFF_X1 \buffer_reg[8][0][2][15]  (.D(\input_filter[0][2] [15]), .CK(n_58_8), 
      .Q(\buffer[8][0][2] [15]), .QN());
   DFF_X1 \buffer_reg[8][0][2][14]  (.D(\input_filter[0][2] [14]), .CK(n_58_8), 
      .Q(\buffer[8][0][2] [14]), .QN());
   DFF_X1 \buffer_reg[8][0][2][13]  (.D(\input_filter[0][2] [13]), .CK(n_58_8), 
      .Q(\buffer[8][0][2] [13]), .QN());
   DFF_X1 \buffer_reg[8][0][2][12]  (.D(\input_filter[0][2] [12]), .CK(n_58_8), 
      .Q(\buffer[8][0][2] [12]), .QN());
   DFF_X1 \buffer_reg[8][0][2][11]  (.D(\input_filter[0][2] [11]), .CK(n_58_8), 
      .Q(\buffer[8][0][2] [11]), .QN());
   DFF_X1 \buffer_reg[8][0][2][10]  (.D(\input_filter[0][2] [10]), .CK(n_58_8), 
      .Q(\buffer[8][0][2] [10]), .QN());
   DFF_X1 \buffer_reg[8][0][2][9]  (.D(\input_filter[0][2] [9]), .CK(n_58_8), 
      .Q(\buffer[8][0][2] [9]), .QN());
   DFF_X1 \buffer_reg[8][0][2][8]  (.D(\input_filter[0][2] [8]), .CK(n_58_8), 
      .Q(\buffer[8][0][2] [8]), .QN());
   DFF_X1 \buffer_reg[8][0][2][7]  (.D(\input_filter[0][2] [7]), .CK(n_58_8), 
      .Q(\buffer[8][0][2] [7]), .QN());
   DFF_X1 \buffer_reg[8][0][2][6]  (.D(\input_filter[0][2] [6]), .CK(n_58_8), 
      .Q(\buffer[8][0][2] [6]), .QN());
   DFF_X1 \buffer_reg[8][0][2][5]  (.D(\input_filter[0][2] [5]), .CK(n_58_8), 
      .Q(\buffer[8][0][2] [5]), .QN());
   DFF_X1 \buffer_reg[8][0][2][4]  (.D(\input_filter[0][2] [4]), .CK(n_58_8), 
      .Q(\buffer[8][0][2] [4]), .QN());
   DFF_X1 \buffer_reg[8][0][2][3]  (.D(\input_filter[0][2] [3]), .CK(n_58_8), 
      .Q(\buffer[8][0][2] [3]), .QN());
   DFF_X1 \buffer_reg[8][0][2][2]  (.D(\input_filter[0][2] [2]), .CK(n_58_8), 
      .Q(\buffer[8][0][2] [2]), .QN());
   DFF_X1 \buffer_reg[8][0][2][1]  (.D(\input_filter[0][2] [1]), .CK(n_58_8), 
      .Q(\buffer[8][0][2] [1]), .QN());
   DFF_X1 \buffer_reg[8][0][2][0]  (.D(\input_filter[0][2] [0]), .CK(n_58_8), 
      .Q(\buffer[8][0][2] [0]), .QN());
   DFF_X1 \buffer_reg[7][0][2][15]  (.D(\input_filter[0][2] [15]), .CK(n_58_7), 
      .Q(\buffer[7][0][2] [15]), .QN());
   DFF_X1 \buffer_reg[7][0][2][14]  (.D(\input_filter[0][2] [14]), .CK(n_58_7), 
      .Q(\buffer[7][0][2] [14]), .QN());
   DFF_X1 \buffer_reg[7][0][2][13]  (.D(\input_filter[0][2] [13]), .CK(n_58_7), 
      .Q(\buffer[7][0][2] [13]), .QN());
   DFF_X1 \buffer_reg[7][0][2][12]  (.D(\input_filter[0][2] [12]), .CK(n_58_7), 
      .Q(\buffer[7][0][2] [12]), .QN());
   DFF_X1 \buffer_reg[7][0][2][11]  (.D(\input_filter[0][2] [11]), .CK(n_58_7), 
      .Q(\buffer[7][0][2] [11]), .QN());
   DFF_X1 \buffer_reg[7][0][2][10]  (.D(\input_filter[0][2] [10]), .CK(n_58_7), 
      .Q(\buffer[7][0][2] [10]), .QN());
   DFF_X1 \buffer_reg[7][0][2][9]  (.D(\input_filter[0][2] [9]), .CK(n_58_7), 
      .Q(\buffer[7][0][2] [9]), .QN());
   DFF_X1 \buffer_reg[7][0][2][8]  (.D(\input_filter[0][2] [8]), .CK(n_58_7), 
      .Q(\buffer[7][0][2] [8]), .QN());
   DFF_X1 \buffer_reg[7][0][2][7]  (.D(\input_filter[0][2] [7]), .CK(n_58_7), 
      .Q(\buffer[7][0][2] [7]), .QN());
   DFF_X1 \buffer_reg[7][0][2][6]  (.D(\input_filter[0][2] [6]), .CK(n_58_7), 
      .Q(\buffer[7][0][2] [6]), .QN());
   DFF_X1 \buffer_reg[7][0][2][5]  (.D(\input_filter[0][2] [5]), .CK(n_58_7), 
      .Q(\buffer[7][0][2] [5]), .QN());
   DFF_X1 \buffer_reg[7][0][2][4]  (.D(\input_filter[0][2] [4]), .CK(n_58_7), 
      .Q(\buffer[7][0][2] [4]), .QN());
   DFF_X1 \buffer_reg[7][0][2][3]  (.D(\input_filter[0][2] [3]), .CK(n_58_7), 
      .Q(\buffer[7][0][2] [3]), .QN());
   DFF_X1 \buffer_reg[7][0][2][2]  (.D(\input_filter[0][2] [2]), .CK(n_58_7), 
      .Q(\buffer[7][0][2] [2]), .QN());
   DFF_X1 \buffer_reg[7][0][2][1]  (.D(\input_filter[0][2] [1]), .CK(n_58_7), 
      .Q(\buffer[7][0][2] [1]), .QN());
   DFF_X1 \buffer_reg[7][0][2][0]  (.D(\input_filter[0][2] [0]), .CK(n_58_7), 
      .Q(\buffer[7][0][2] [0]), .QN());
   DFF_X1 \buffer_reg[0][0][2][15]  (.D(\input_filter[0][2] [15]), .CK(n_58_0), 
      .Q(\buffer[0][0][2] [15]), .QN());
   DFF_X1 \buffer_reg[0][0][2][14]  (.D(\input_filter[0][2] [14]), .CK(n_58_0), 
      .Q(\buffer[0][0][2] [14]), .QN());
   DFF_X1 \buffer_reg[0][0][2][13]  (.D(\input_filter[0][2] [13]), .CK(n_58_0), 
      .Q(\buffer[0][0][2] [13]), .QN());
   DFF_X1 \buffer_reg[0][0][2][12]  (.D(\input_filter[0][2] [12]), .CK(n_58_0), 
      .Q(\buffer[0][0][2] [12]), .QN());
   DFF_X1 \buffer_reg[0][0][2][11]  (.D(\input_filter[0][2] [11]), .CK(n_58_0), 
      .Q(\buffer[0][0][2] [11]), .QN());
   DFF_X1 \buffer_reg[0][0][2][10]  (.D(\input_filter[0][2] [10]), .CK(n_58_0), 
      .Q(\buffer[0][0][2] [10]), .QN());
   DFF_X1 \buffer_reg[0][0][2][9]  (.D(\input_filter[0][2] [9]), .CK(n_58_0), 
      .Q(\buffer[0][0][2] [9]), .QN());
   DFF_X1 \buffer_reg[0][0][2][8]  (.D(\input_filter[0][2] [8]), .CK(n_58_0), 
      .Q(\buffer[0][0][2] [8]), .QN());
   DFF_X1 \buffer_reg[0][0][2][7]  (.D(\input_filter[0][2] [7]), .CK(n_58_0), 
      .Q(\buffer[0][0][2] [7]), .QN());
   DFF_X1 \buffer_reg[0][0][2][6]  (.D(\input_filter[0][2] [6]), .CK(n_58_0), 
      .Q(\buffer[0][0][2] [6]), .QN());
   DFF_X1 \buffer_reg[0][0][2][5]  (.D(\input_filter[0][2] [5]), .CK(n_58_0), 
      .Q(\buffer[0][0][2] [5]), .QN());
   DFF_X1 \buffer_reg[0][0][2][4]  (.D(\input_filter[0][2] [4]), .CK(n_58_0), 
      .Q(\buffer[0][0][2] [4]), .QN());
   DFF_X1 \buffer_reg[0][0][2][3]  (.D(\input_filter[0][2] [3]), .CK(n_58_0), 
      .Q(\buffer[0][0][2] [3]), .QN());
   DFF_X1 \buffer_reg[0][0][2][2]  (.D(\input_filter[0][2] [2]), .CK(n_58_0), 
      .Q(\buffer[0][0][2] [2]), .QN());
   DFF_X1 \buffer_reg[0][0][2][1]  (.D(\input_filter[0][2] [1]), .CK(n_58_0), 
      .Q(\buffer[0][0][2] [1]), .QN());
   DFF_X1 \buffer_reg[0][0][2][0]  (.D(\input_filter[0][2] [0]), .CK(n_58_0), 
      .Q(\buffer[0][0][2] [0]), .QN());
   CLKGATETST_X1 \clk_gate_buffer_reg[0][1][3]_reg  (.CK(read), .E(n_0), 
      .SE(1'b0), .GCK(n_58_0));
   CLKGATETST_X1 \clk_gate_buffer_reg[1][1][3]_reg  (.CK(read), .E(n_1), 
      .SE(1'b0), .GCK(n_58_1));
   CLKGATETST_X1 \clk_gate_buffer_reg[2][1][3]_reg  (.CK(read), .E(n_2), 
      .SE(1'b0), .GCK(n_58_2));
   CLKGATETST_X1 \clk_gate_buffer_reg[3][1][3]_reg  (.CK(read), .E(n_3), 
      .SE(1'b0), .GCK(n_58_3));
   CLKGATETST_X1 \clk_gate_buffer_reg[4][1][3]_reg  (.CK(read), .E(n_4), 
      .SE(1'b0), .GCK(n_58_4));
   CLKGATETST_X1 \clk_gate_buffer_reg[5][1][3]_reg  (.CK(read), .E(n_5), 
      .SE(1'b0), .GCK(n_58_5));
   CLKGATETST_X1 \clk_gate_buffer_reg[7][1][3]_reg  (.CK(read), .E(n_7), 
      .SE(1'b0), .GCK(n_58_7));
   CLKGATETST_X1 \clk_gate_buffer_reg[8][1][3]_reg  (.CK(read), .E(n_8), 
      .SE(1'b0), .GCK(n_58_8));
   CLKGATETST_X1 \clk_gate_buffer_reg[9][1][3]_reg  (.CK(read), .E(n_9), 
      .SE(1'b0), .GCK(n_58_9));
   CLKGATETST_X1 \clk_gate_buffer_reg[10][1][3]_reg  (.CK(read), .E(n_10), 
      .SE(1'b0), .GCK(n_58_10));
   CLKGATETST_X1 \clk_gate_buffer_reg[11][1][3]_reg  (.CK(read), .E(n_11), 
      .SE(1'b0), .GCK(n_58_11));
   CLKGATETST_X1 \clk_gate_buffer_reg[12][1][3]_reg  (.CK(read), .E(n_12), 
      .SE(1'b0), .GCK(n_58_12));
   CLKGATETST_X1 \clk_gate_buffer_reg[13][1][3]_reg  (.CK(read), .E(n_13), 
      .SE(1'b0), .GCK(n_58_13));
   CLKGATETST_X1 \clk_gate_buffer_reg[14][1][3]_reg  (.CK(read), .E(n_14), 
      .SE(1'b0), .GCK(n_58_14));
   DFF_X1 \buffer_reg[0][1][4][15]  (.D(\input_filter[1][4] [15]), .CK(n_59_0), 
      .Q(\buffer[0][1][4] [15]), .QN());
   DFF_X1 \buffer_reg[0][1][4][14]  (.D(\input_filter[1][4] [14]), .CK(n_59_0), 
      .Q(\buffer[0][1][4] [14]), .QN());
   DFF_X1 \buffer_reg[0][1][4][13]  (.D(\input_filter[1][4] [13]), .CK(n_59_0), 
      .Q(\buffer[0][1][4] [13]), .QN());
   DFF_X1 \buffer_reg[0][1][4][12]  (.D(\input_filter[1][4] [12]), .CK(n_59_0), 
      .Q(\buffer[0][1][4] [12]), .QN());
   DFF_X1 \buffer_reg[0][1][4][11]  (.D(\input_filter[1][4] [11]), .CK(n_59_0), 
      .Q(\buffer[0][1][4] [11]), .QN());
   DFF_X1 \buffer_reg[0][1][4][10]  (.D(\input_filter[1][4] [10]), .CK(n_59_0), 
      .Q(\buffer[0][1][4] [10]), .QN());
   DFF_X1 \buffer_reg[0][1][4][9]  (.D(\input_filter[1][4] [9]), .CK(n_59_0), 
      .Q(\buffer[0][1][4] [9]), .QN());
   DFF_X1 \buffer_reg[0][1][4][8]  (.D(\input_filter[1][4] [8]), .CK(n_59_0), 
      .Q(\buffer[0][1][4] [8]), .QN());
   DFF_X1 \buffer_reg[0][1][4][7]  (.D(\input_filter[1][4] [7]), .CK(n_59_0), 
      .Q(\buffer[0][1][4] [7]), .QN());
   DFF_X1 \buffer_reg[0][1][4][6]  (.D(\input_filter[1][4] [6]), .CK(n_59_0), 
      .Q(\buffer[0][1][4] [6]), .QN());
   DFF_X1 \buffer_reg[0][1][4][5]  (.D(\input_filter[1][4] [5]), .CK(n_59_0), 
      .Q(\buffer[0][1][4] [5]), .QN());
   DFF_X1 \buffer_reg[0][1][4][4]  (.D(\input_filter[1][4] [4]), .CK(n_59_0), 
      .Q(\buffer[0][1][4] [4]), .QN());
   DFF_X1 \buffer_reg[0][1][4][3]  (.D(\input_filter[1][4] [3]), .CK(n_59_0), 
      .Q(\buffer[0][1][4] [3]), .QN());
   DFF_X1 \buffer_reg[0][1][4][2]  (.D(\input_filter[1][4] [2]), .CK(n_59_0), 
      .Q(\buffer[0][1][4] [2]), .QN());
   DFF_X1 \buffer_reg[0][1][4][1]  (.D(\input_filter[1][4] [1]), .CK(n_59_0), 
      .Q(\buffer[0][1][4] [1]), .QN());
   DFF_X1 \buffer_reg[0][1][4][0]  (.D(\input_filter[1][4] [0]), .CK(n_59_0), 
      .Q(\buffer[0][1][4] [0]), .QN());
   DFF_X1 \buffer_reg[11][1][4][15]  (.D(\input_filter[1][4] [15]), .CK(n_59_1), 
      .Q(\buffer[11][1][4] [15]), .QN());
   DFF_X1 \buffer_reg[11][1][4][14]  (.D(\input_filter[1][4] [14]), .CK(n_59_1), 
      .Q(\buffer[11][1][4] [14]), .QN());
   DFF_X1 \buffer_reg[11][1][4][13]  (.D(\input_filter[1][4] [13]), .CK(n_59_1), 
      .Q(\buffer[11][1][4] [13]), .QN());
   DFF_X1 \buffer_reg[11][1][4][12]  (.D(\input_filter[1][4] [12]), .CK(n_59_1), 
      .Q(\buffer[11][1][4] [12]), .QN());
   DFF_X1 \buffer_reg[11][1][4][11]  (.D(\input_filter[1][4] [11]), .CK(n_59_1), 
      .Q(\buffer[11][1][4] [11]), .QN());
   DFF_X1 \buffer_reg[11][1][4][10]  (.D(\input_filter[1][4] [10]), .CK(n_59_1), 
      .Q(\buffer[11][1][4] [10]), .QN());
   DFF_X1 \buffer_reg[11][1][4][9]  (.D(\input_filter[1][4] [9]), .CK(n_59_1), 
      .Q(\buffer[11][1][4] [9]), .QN());
   DFF_X1 \buffer_reg[11][1][4][8]  (.D(\input_filter[1][4] [8]), .CK(n_59_1), 
      .Q(\buffer[11][1][4] [8]), .QN());
   DFF_X1 \buffer_reg[11][1][4][7]  (.D(\input_filter[1][4] [7]), .CK(n_59_1), 
      .Q(\buffer[11][1][4] [7]), .QN());
   DFF_X1 \buffer_reg[11][1][4][6]  (.D(\input_filter[1][4] [6]), .CK(n_59_1), 
      .Q(\buffer[11][1][4] [6]), .QN());
   DFF_X1 \buffer_reg[11][1][4][5]  (.D(\input_filter[1][4] [5]), .CK(n_59_1), 
      .Q(\buffer[11][1][4] [5]), .QN());
   DFF_X1 \buffer_reg[11][1][4][4]  (.D(\input_filter[1][4] [4]), .CK(n_59_1), 
      .Q(\buffer[11][1][4] [4]), .QN());
   DFF_X1 \buffer_reg[11][1][4][3]  (.D(\input_filter[1][4] [3]), .CK(n_59_1), 
      .Q(\buffer[11][1][4] [3]), .QN());
   DFF_X1 \buffer_reg[11][1][4][2]  (.D(\input_filter[1][4] [2]), .CK(n_59_1), 
      .Q(\buffer[11][1][4] [2]), .QN());
   DFF_X1 \buffer_reg[11][1][4][1]  (.D(\input_filter[1][4] [1]), .CK(n_59_1), 
      .Q(\buffer[11][1][4] [1]), .QN());
   DFF_X1 \buffer_reg[11][1][4][0]  (.D(\input_filter[1][4] [0]), .CK(n_59_1), 
      .Q(\buffer[11][1][4] [0]), .QN());
   DFF_X1 \buffer_reg[12][1][4][15]  (.D(\input_filter[1][4] [15]), .CK(n_59_2), 
      .Q(\buffer[12][1][4] [15]), .QN());
   DFF_X1 \buffer_reg[12][1][4][14]  (.D(\input_filter[1][4] [14]), .CK(n_59_2), 
      .Q(\buffer[12][1][4] [14]), .QN());
   DFF_X1 \buffer_reg[12][1][4][13]  (.D(\input_filter[1][4] [13]), .CK(n_59_2), 
      .Q(\buffer[12][1][4] [13]), .QN());
   DFF_X1 \buffer_reg[12][1][4][12]  (.D(\input_filter[1][4] [12]), .CK(n_59_2), 
      .Q(\buffer[12][1][4] [12]), .QN());
   DFF_X1 \buffer_reg[12][1][4][11]  (.D(\input_filter[1][4] [11]), .CK(n_59_2), 
      .Q(\buffer[12][1][4] [11]), .QN());
   DFF_X1 \buffer_reg[12][1][4][10]  (.D(\input_filter[1][4] [10]), .CK(n_59_2), 
      .Q(\buffer[12][1][4] [10]), .QN());
   DFF_X1 \buffer_reg[12][1][4][9]  (.D(\input_filter[1][4] [9]), .CK(n_59_2), 
      .Q(\buffer[12][1][4] [9]), .QN());
   DFF_X1 \buffer_reg[12][1][4][8]  (.D(\input_filter[1][4] [8]), .CK(n_59_2), 
      .Q(\buffer[12][1][4] [8]), .QN());
   DFF_X1 \buffer_reg[12][1][4][7]  (.D(\input_filter[1][4] [7]), .CK(n_59_2), 
      .Q(\buffer[12][1][4] [7]), .QN());
   DFF_X1 \buffer_reg[12][1][4][6]  (.D(\input_filter[1][4] [6]), .CK(n_59_2), 
      .Q(\buffer[12][1][4] [6]), .QN());
   DFF_X1 \buffer_reg[12][1][4][5]  (.D(\input_filter[1][4] [5]), .CK(n_59_2), 
      .Q(\buffer[12][1][4] [5]), .QN());
   DFF_X1 \buffer_reg[12][1][4][4]  (.D(\input_filter[1][4] [4]), .CK(n_59_2), 
      .Q(\buffer[12][1][4] [4]), .QN());
   DFF_X1 \buffer_reg[12][1][4][3]  (.D(\input_filter[1][4] [3]), .CK(n_59_2), 
      .Q(\buffer[12][1][4] [3]), .QN());
   DFF_X1 \buffer_reg[12][1][4][2]  (.D(\input_filter[1][4] [2]), .CK(n_59_2), 
      .Q(\buffer[12][1][4] [2]), .QN());
   DFF_X1 \buffer_reg[12][1][4][1]  (.D(\input_filter[1][4] [1]), .CK(n_59_2), 
      .Q(\buffer[12][1][4] [1]), .QN());
   DFF_X1 \buffer_reg[12][1][4][0]  (.D(\input_filter[1][4] [0]), .CK(n_59_2), 
      .Q(\buffer[12][1][4] [0]), .QN());
   DFF_X1 \buffer_reg[13][1][4][15]  (.D(\input_filter[1][4] [15]), .CK(n_59_3), 
      .Q(\buffer[13][1][4] [15]), .QN());
   DFF_X1 \buffer_reg[13][1][4][14]  (.D(\input_filter[1][4] [14]), .CK(n_59_3), 
      .Q(\buffer[13][1][4] [14]), .QN());
   DFF_X1 \buffer_reg[13][1][4][13]  (.D(\input_filter[1][4] [13]), .CK(n_59_3), 
      .Q(\buffer[13][1][4] [13]), .QN());
   DFF_X1 \buffer_reg[13][1][4][12]  (.D(\input_filter[1][4] [12]), .CK(n_59_3), 
      .Q(\buffer[13][1][4] [12]), .QN());
   DFF_X1 \buffer_reg[13][1][4][11]  (.D(\input_filter[1][4] [11]), .CK(n_59_3), 
      .Q(\buffer[13][1][4] [11]), .QN());
   DFF_X1 \buffer_reg[13][1][4][10]  (.D(\input_filter[1][4] [10]), .CK(n_59_3), 
      .Q(\buffer[13][1][4] [10]), .QN());
   DFF_X1 \buffer_reg[13][1][4][9]  (.D(\input_filter[1][4] [9]), .CK(n_59_3), 
      .Q(\buffer[13][1][4] [9]), .QN());
   DFF_X1 \buffer_reg[13][1][4][8]  (.D(\input_filter[1][4] [8]), .CK(n_59_3), 
      .Q(\buffer[13][1][4] [8]), .QN());
   DFF_X1 \buffer_reg[13][1][4][7]  (.D(\input_filter[1][4] [7]), .CK(n_59_3), 
      .Q(\buffer[13][1][4] [7]), .QN());
   DFF_X1 \buffer_reg[13][1][4][6]  (.D(\input_filter[1][4] [6]), .CK(n_59_3), 
      .Q(\buffer[13][1][4] [6]), .QN());
   DFF_X1 \buffer_reg[13][1][4][5]  (.D(\input_filter[1][4] [5]), .CK(n_59_3), 
      .Q(\buffer[13][1][4] [5]), .QN());
   DFF_X1 \buffer_reg[13][1][4][4]  (.D(\input_filter[1][4] [4]), .CK(n_59_3), 
      .Q(\buffer[13][1][4] [4]), .QN());
   DFF_X1 \buffer_reg[13][1][4][3]  (.D(\input_filter[1][4] [3]), .CK(n_59_3), 
      .Q(\buffer[13][1][4] [3]), .QN());
   DFF_X1 \buffer_reg[13][1][4][2]  (.D(\input_filter[1][4] [2]), .CK(n_59_3), 
      .Q(\buffer[13][1][4] [2]), .QN());
   DFF_X1 \buffer_reg[13][1][4][1]  (.D(\input_filter[1][4] [1]), .CK(n_59_3), 
      .Q(\buffer[13][1][4] [1]), .QN());
   DFF_X1 \buffer_reg[13][1][4][0]  (.D(\input_filter[1][4] [0]), .CK(n_59_3), 
      .Q(\buffer[13][1][4] [0]), .QN());
   DFF_X1 \buffer_reg[14][1][4][15]  (.D(\input_filter[1][4] [15]), .CK(n_59_4), 
      .Q(\buffer[14][1][4] [15]), .QN());
   DFF_X1 \buffer_reg[14][1][4][14]  (.D(\input_filter[1][4] [14]), .CK(n_59_4), 
      .Q(\buffer[14][1][4] [14]), .QN());
   DFF_X1 \buffer_reg[14][1][4][13]  (.D(\input_filter[1][4] [13]), .CK(n_59_4), 
      .Q(\buffer[14][1][4] [13]), .QN());
   DFF_X1 \buffer_reg[14][1][4][12]  (.D(\input_filter[1][4] [12]), .CK(n_59_4), 
      .Q(\buffer[14][1][4] [12]), .QN());
   DFF_X1 \buffer_reg[14][1][4][11]  (.D(\input_filter[1][4] [11]), .CK(n_59_4), 
      .Q(\buffer[14][1][4] [11]), .QN());
   DFF_X1 \buffer_reg[14][1][4][10]  (.D(\input_filter[1][4] [10]), .CK(n_59_4), 
      .Q(\buffer[14][1][4] [10]), .QN());
   DFF_X1 \buffer_reg[14][1][4][9]  (.D(\input_filter[1][4] [9]), .CK(n_59_4), 
      .Q(\buffer[14][1][4] [9]), .QN());
   DFF_X1 \buffer_reg[14][1][4][8]  (.D(\input_filter[1][4] [8]), .CK(n_59_4), 
      .Q(\buffer[14][1][4] [8]), .QN());
   DFF_X1 \buffer_reg[14][1][4][7]  (.D(\input_filter[1][4] [7]), .CK(n_59_4), 
      .Q(\buffer[14][1][4] [7]), .QN());
   DFF_X1 \buffer_reg[14][1][4][6]  (.D(\input_filter[1][4] [6]), .CK(n_59_4), 
      .Q(\buffer[14][1][4] [6]), .QN());
   DFF_X1 \buffer_reg[14][1][4][5]  (.D(\input_filter[1][4] [5]), .CK(n_59_4), 
      .Q(\buffer[14][1][4] [5]), .QN());
   DFF_X1 \buffer_reg[14][1][4][4]  (.D(\input_filter[1][4] [4]), .CK(n_59_4), 
      .Q(\buffer[14][1][4] [4]), .QN());
   DFF_X1 \buffer_reg[14][1][4][3]  (.D(\input_filter[1][4] [3]), .CK(n_59_4), 
      .Q(\buffer[14][1][4] [3]), .QN());
   DFF_X1 \buffer_reg[14][1][4][2]  (.D(\input_filter[1][4] [2]), .CK(n_59_4), 
      .Q(\buffer[14][1][4] [2]), .QN());
   DFF_X1 \buffer_reg[14][1][4][1]  (.D(\input_filter[1][4] [1]), .CK(n_59_4), 
      .Q(\buffer[14][1][4] [1]), .QN());
   DFF_X1 \buffer_reg[14][1][4][0]  (.D(\input_filter[1][4] [0]), .CK(n_59_4), 
      .Q(\buffer[14][1][4] [0]), .QN());
   DFF_X1 \buffer_reg[15][1][4][15]  (.D(\input_filter[1][4] [15]), .CK(n_59_5), 
      .Q(\buffer[15][1][4] [15]), .QN());
   DFF_X1 \buffer_reg[15][1][4][14]  (.D(\input_filter[1][4] [14]), .CK(n_59_5), 
      .Q(\buffer[15][1][4] [14]), .QN());
   DFF_X1 \buffer_reg[15][1][4][13]  (.D(\input_filter[1][4] [13]), .CK(n_59_5), 
      .Q(\buffer[15][1][4] [13]), .QN());
   DFF_X1 \buffer_reg[15][1][4][12]  (.D(\input_filter[1][4] [12]), .CK(n_59_5), 
      .Q(\buffer[15][1][4] [12]), .QN());
   DFF_X1 \buffer_reg[15][1][4][11]  (.D(\input_filter[1][4] [11]), .CK(n_59_5), 
      .Q(\buffer[15][1][4] [11]), .QN());
   DFF_X1 \buffer_reg[15][1][4][10]  (.D(\input_filter[1][4] [10]), .CK(n_59_5), 
      .Q(\buffer[15][1][4] [10]), .QN());
   DFF_X1 \buffer_reg[15][1][4][9]  (.D(\input_filter[1][4] [9]), .CK(n_59_5), 
      .Q(\buffer[15][1][4] [9]), .QN());
   DFF_X1 \buffer_reg[15][1][4][8]  (.D(\input_filter[1][4] [8]), .CK(n_59_5), 
      .Q(\buffer[15][1][4] [8]), .QN());
   DFF_X1 \buffer_reg[15][1][4][7]  (.D(\input_filter[1][4] [7]), .CK(n_59_5), 
      .Q(\buffer[15][1][4] [7]), .QN());
   DFF_X1 \buffer_reg[15][1][4][6]  (.D(\input_filter[1][4] [6]), .CK(n_59_5), 
      .Q(\buffer[15][1][4] [6]), .QN());
   DFF_X1 \buffer_reg[15][1][4][5]  (.D(\input_filter[1][4] [5]), .CK(n_59_5), 
      .Q(\buffer[15][1][4] [5]), .QN());
   DFF_X1 \buffer_reg[15][1][4][4]  (.D(\input_filter[1][4] [4]), .CK(n_59_5), 
      .Q(\buffer[15][1][4] [4]), .QN());
   DFF_X1 \buffer_reg[15][1][4][3]  (.D(\input_filter[1][4] [3]), .CK(n_59_5), 
      .Q(\buffer[15][1][4] [3]), .QN());
   DFF_X1 \buffer_reg[15][1][4][2]  (.D(\input_filter[1][4] [2]), .CK(n_59_5), 
      .Q(\buffer[15][1][4] [2]), .QN());
   DFF_X1 \buffer_reg[15][1][4][1]  (.D(\input_filter[1][4] [1]), .CK(n_59_5), 
      .Q(\buffer[15][1][4] [1]), .QN());
   DFF_X1 \buffer_reg[15][1][4][0]  (.D(\input_filter[1][4] [0]), .CK(n_59_5), 
      .Q(\buffer[15][1][4] [0]), .QN());
   DFF_X1 \buffer_reg[0][2][0][15]  (.D(\input_filter[2][0] [15]), .CK(n_59_0), 
      .Q(\buffer[0][2][0] [15]), .QN());
   DFF_X1 \buffer_reg[0][2][0][14]  (.D(\input_filter[2][0] [14]), .CK(n_59_0), 
      .Q(\buffer[0][2][0] [14]), .QN());
   DFF_X1 \buffer_reg[0][2][0][13]  (.D(\input_filter[2][0] [13]), .CK(n_59_0), 
      .Q(\buffer[0][2][0] [13]), .QN());
   DFF_X1 \buffer_reg[0][2][0][12]  (.D(\input_filter[2][0] [12]), .CK(n_59_0), 
      .Q(\buffer[0][2][0] [12]), .QN());
   DFF_X1 \buffer_reg[0][2][0][11]  (.D(\input_filter[2][0] [11]), .CK(n_59_0), 
      .Q(\buffer[0][2][0] [11]), .QN());
   DFF_X1 \buffer_reg[0][2][0][10]  (.D(\input_filter[2][0] [10]), .CK(n_59_0), 
      .Q(\buffer[0][2][0] [10]), .QN());
   DFF_X1 \buffer_reg[0][2][0][9]  (.D(\input_filter[2][0] [9]), .CK(n_59_0), 
      .Q(\buffer[0][2][0] [9]), .QN());
   DFF_X1 \buffer_reg[0][2][0][8]  (.D(\input_filter[2][0] [8]), .CK(n_59_0), 
      .Q(\buffer[0][2][0] [8]), .QN());
   DFF_X1 \buffer_reg[0][2][0][7]  (.D(\input_filter[2][0] [7]), .CK(n_59_0), 
      .Q(\buffer[0][2][0] [7]), .QN());
   DFF_X1 \buffer_reg[0][2][0][6]  (.D(\input_filter[2][0] [6]), .CK(n_59_0), 
      .Q(\buffer[0][2][0] [6]), .QN());
   DFF_X1 \buffer_reg[0][2][0][5]  (.D(\input_filter[2][0] [5]), .CK(n_59_0), 
      .Q(\buffer[0][2][0] [5]), .QN());
   DFF_X1 \buffer_reg[0][2][0][4]  (.D(\input_filter[2][0] [4]), .CK(n_59_0), 
      .Q(\buffer[0][2][0] [4]), .QN());
   DFF_X1 \buffer_reg[0][2][0][3]  (.D(\input_filter[2][0] [3]), .CK(n_59_0), 
      .Q(\buffer[0][2][0] [3]), .QN());
   DFF_X1 \buffer_reg[0][2][0][2]  (.D(\input_filter[2][0] [2]), .CK(n_59_0), 
      .Q(\buffer[0][2][0] [2]), .QN());
   DFF_X1 \buffer_reg[0][2][0][1]  (.D(\input_filter[2][0] [1]), .CK(n_59_0), 
      .Q(\buffer[0][2][0] [1]), .QN());
   DFF_X1 \buffer_reg[0][2][0][0]  (.D(\input_filter[2][0] [0]), .CK(n_59_0), 
      .Q(\buffer[0][2][0] [0]), .QN());
   DFF_X1 \buffer_reg[1][2][0][15]  (.D(\input_filter[2][0] [15]), .CK(n_59_7), 
      .Q(\buffer[1][2][0] [15]), .QN());
   DFF_X1 \buffer_reg[1][2][0][14]  (.D(\input_filter[2][0] [14]), .CK(n_59_7), 
      .Q(\buffer[1][2][0] [14]), .QN());
   DFF_X1 \buffer_reg[1][2][0][13]  (.D(\input_filter[2][0] [13]), .CK(n_59_7), 
      .Q(\buffer[1][2][0] [13]), .QN());
   DFF_X1 \buffer_reg[1][2][0][12]  (.D(\input_filter[2][0] [12]), .CK(n_59_7), 
      .Q(\buffer[1][2][0] [12]), .QN());
   DFF_X1 \buffer_reg[1][2][0][11]  (.D(\input_filter[2][0] [11]), .CK(n_59_7), 
      .Q(\buffer[1][2][0] [11]), .QN());
   DFF_X1 \buffer_reg[1][2][0][10]  (.D(\input_filter[2][0] [10]), .CK(n_59_7), 
      .Q(\buffer[1][2][0] [10]), .QN());
   DFF_X1 \buffer_reg[1][2][0][9]  (.D(\input_filter[2][0] [9]), .CK(n_59_7), 
      .Q(\buffer[1][2][0] [9]), .QN());
   DFF_X1 \buffer_reg[1][2][0][8]  (.D(\input_filter[2][0] [8]), .CK(n_59_7), 
      .Q(\buffer[1][2][0] [8]), .QN());
   DFF_X1 \buffer_reg[1][2][0][7]  (.D(\input_filter[2][0] [7]), .CK(n_59_7), 
      .Q(\buffer[1][2][0] [7]), .QN());
   DFF_X1 \buffer_reg[1][2][0][6]  (.D(\input_filter[2][0] [6]), .CK(n_59_7), 
      .Q(\buffer[1][2][0] [6]), .QN());
   DFF_X1 \buffer_reg[1][2][0][5]  (.D(\input_filter[2][0] [5]), .CK(n_59_7), 
      .Q(\buffer[1][2][0] [5]), .QN());
   DFF_X1 \buffer_reg[1][2][0][4]  (.D(\input_filter[2][0] [4]), .CK(n_59_7), 
      .Q(\buffer[1][2][0] [4]), .QN());
   DFF_X1 \buffer_reg[1][2][0][3]  (.D(\input_filter[2][0] [3]), .CK(n_59_7), 
      .Q(\buffer[1][2][0] [3]), .QN());
   DFF_X1 \buffer_reg[1][2][0][2]  (.D(\input_filter[2][0] [2]), .CK(n_59_7), 
      .Q(\buffer[1][2][0] [2]), .QN());
   DFF_X1 \buffer_reg[1][2][0][1]  (.D(\input_filter[2][0] [1]), .CK(n_59_7), 
      .Q(\buffer[1][2][0] [1]), .QN());
   DFF_X1 \buffer_reg[1][2][0][0]  (.D(\input_filter[2][0] [0]), .CK(n_59_7), 
      .Q(\buffer[1][2][0] [0]), .QN());
   DFF_X1 \buffer_reg[2][2][0][15]  (.D(\input_filter[2][0] [15]), .CK(n_59_8), 
      .Q(\buffer[2][2][0] [15]), .QN());
   DFF_X1 \buffer_reg[2][2][0][14]  (.D(\input_filter[2][0] [14]), .CK(n_59_8), 
      .Q(\buffer[2][2][0] [14]), .QN());
   DFF_X1 \buffer_reg[2][2][0][13]  (.D(\input_filter[2][0] [13]), .CK(n_59_8), 
      .Q(\buffer[2][2][0] [13]), .QN());
   DFF_X1 \buffer_reg[2][2][0][12]  (.D(\input_filter[2][0] [12]), .CK(n_59_8), 
      .Q(\buffer[2][2][0] [12]), .QN());
   DFF_X1 \buffer_reg[2][2][0][11]  (.D(\input_filter[2][0] [11]), .CK(n_59_8), 
      .Q(\buffer[2][2][0] [11]), .QN());
   DFF_X1 \buffer_reg[2][2][0][10]  (.D(\input_filter[2][0] [10]), .CK(n_59_8), 
      .Q(\buffer[2][2][0] [10]), .QN());
   DFF_X1 \buffer_reg[2][2][0][9]  (.D(\input_filter[2][0] [9]), .CK(n_59_8), 
      .Q(\buffer[2][2][0] [9]), .QN());
   DFF_X1 \buffer_reg[2][2][0][8]  (.D(\input_filter[2][0] [8]), .CK(n_59_8), 
      .Q(\buffer[2][2][0] [8]), .QN());
   DFF_X1 \buffer_reg[2][2][0][7]  (.D(\input_filter[2][0] [7]), .CK(n_59_8), 
      .Q(\buffer[2][2][0] [7]), .QN());
   DFF_X1 \buffer_reg[2][2][0][6]  (.D(\input_filter[2][0] [6]), .CK(n_59_8), 
      .Q(\buffer[2][2][0] [6]), .QN());
   DFF_X1 \buffer_reg[2][2][0][5]  (.D(\input_filter[2][0] [5]), .CK(n_59_8), 
      .Q(\buffer[2][2][0] [5]), .QN());
   DFF_X1 \buffer_reg[2][2][0][4]  (.D(\input_filter[2][0] [4]), .CK(n_59_8), 
      .Q(\buffer[2][2][0] [4]), .QN());
   DFF_X1 \buffer_reg[2][2][0][3]  (.D(\input_filter[2][0] [3]), .CK(n_59_8), 
      .Q(\buffer[2][2][0] [3]), .QN());
   DFF_X1 \buffer_reg[2][2][0][2]  (.D(\input_filter[2][0] [2]), .CK(n_59_8), 
      .Q(\buffer[2][2][0] [2]), .QN());
   DFF_X1 \buffer_reg[2][2][0][1]  (.D(\input_filter[2][0] [1]), .CK(n_59_8), 
      .Q(\buffer[2][2][0] [1]), .QN());
   DFF_X1 \buffer_reg[2][2][0][0]  (.D(\input_filter[2][0] [0]), .CK(n_59_8), 
      .Q(\buffer[2][2][0] [0]), .QN());
   DFF_X1 \buffer_reg[3][2][0][15]  (.D(\input_filter[2][0] [15]), .CK(n_59_9), 
      .Q(\buffer[3][2][0] [15]), .QN());
   DFF_X1 \buffer_reg[3][2][0][14]  (.D(\input_filter[2][0] [14]), .CK(n_59_9), 
      .Q(\buffer[3][2][0] [14]), .QN());
   DFF_X1 \buffer_reg[3][2][0][13]  (.D(\input_filter[2][0] [13]), .CK(n_59_9), 
      .Q(\buffer[3][2][0] [13]), .QN());
   DFF_X1 \buffer_reg[3][2][0][12]  (.D(\input_filter[2][0] [12]), .CK(n_59_9), 
      .Q(\buffer[3][2][0] [12]), .QN());
   DFF_X1 \buffer_reg[3][2][0][11]  (.D(\input_filter[2][0] [11]), .CK(n_59_9), 
      .Q(\buffer[3][2][0] [11]), .QN());
   DFF_X1 \buffer_reg[3][2][0][10]  (.D(\input_filter[2][0] [10]), .CK(n_59_9), 
      .Q(\buffer[3][2][0] [10]), .QN());
   DFF_X1 \buffer_reg[3][2][0][9]  (.D(\input_filter[2][0] [9]), .CK(n_59_9), 
      .Q(\buffer[3][2][0] [9]), .QN());
   DFF_X1 \buffer_reg[3][2][0][8]  (.D(\input_filter[2][0] [8]), .CK(n_59_9), 
      .Q(\buffer[3][2][0] [8]), .QN());
   DFF_X1 \buffer_reg[3][2][0][7]  (.D(\input_filter[2][0] [7]), .CK(n_59_9), 
      .Q(\buffer[3][2][0] [7]), .QN());
   DFF_X1 \buffer_reg[3][2][0][6]  (.D(\input_filter[2][0] [6]), .CK(n_59_9), 
      .Q(\buffer[3][2][0] [6]), .QN());
   DFF_X1 \buffer_reg[3][2][0][5]  (.D(\input_filter[2][0] [5]), .CK(n_59_9), 
      .Q(\buffer[3][2][0] [5]), .QN());
   DFF_X1 \buffer_reg[3][2][0][4]  (.D(\input_filter[2][0] [4]), .CK(n_59_9), 
      .Q(\buffer[3][2][0] [4]), .QN());
   DFF_X1 \buffer_reg[3][2][0][3]  (.D(\input_filter[2][0] [3]), .CK(n_59_9), 
      .Q(\buffer[3][2][0] [3]), .QN());
   DFF_X1 \buffer_reg[3][2][0][2]  (.D(\input_filter[2][0] [2]), .CK(n_59_9), 
      .Q(\buffer[3][2][0] [2]), .QN());
   DFF_X1 \buffer_reg[3][2][0][1]  (.D(\input_filter[2][0] [1]), .CK(n_59_9), 
      .Q(\buffer[3][2][0] [1]), .QN());
   DFF_X1 \buffer_reg[3][2][0][0]  (.D(\input_filter[2][0] [0]), .CK(n_59_9), 
      .Q(\buffer[3][2][0] [0]), .QN());
   DFF_X1 \buffer_reg[4][2][0][15]  (.D(\input_filter[2][0] [15]), .CK(n_59_10), 
      .Q(\buffer[4][2][0] [15]), .QN());
   DFF_X1 \buffer_reg[4][2][0][14]  (.D(\input_filter[2][0] [14]), .CK(n_59_10), 
      .Q(\buffer[4][2][0] [14]), .QN());
   DFF_X1 \buffer_reg[4][2][0][13]  (.D(\input_filter[2][0] [13]), .CK(n_59_10), 
      .Q(\buffer[4][2][0] [13]), .QN());
   DFF_X1 \buffer_reg[4][2][0][12]  (.D(\input_filter[2][0] [12]), .CK(n_59_10), 
      .Q(\buffer[4][2][0] [12]), .QN());
   DFF_X1 \buffer_reg[4][2][0][11]  (.D(\input_filter[2][0] [11]), .CK(n_59_10), 
      .Q(\buffer[4][2][0] [11]), .QN());
   DFF_X1 \buffer_reg[4][2][0][10]  (.D(\input_filter[2][0] [10]), .CK(n_59_10), 
      .Q(\buffer[4][2][0] [10]), .QN());
   DFF_X1 \buffer_reg[4][2][0][9]  (.D(\input_filter[2][0] [9]), .CK(n_59_10), 
      .Q(\buffer[4][2][0] [9]), .QN());
   DFF_X1 \buffer_reg[4][2][0][8]  (.D(\input_filter[2][0] [8]), .CK(n_59_10), 
      .Q(\buffer[4][2][0] [8]), .QN());
   DFF_X1 \buffer_reg[4][2][0][7]  (.D(\input_filter[2][0] [7]), .CK(n_59_10), 
      .Q(\buffer[4][2][0] [7]), .QN());
   DFF_X1 \buffer_reg[4][2][0][6]  (.D(\input_filter[2][0] [6]), .CK(n_59_10), 
      .Q(\buffer[4][2][0] [6]), .QN());
   DFF_X1 \buffer_reg[4][2][0][5]  (.D(\input_filter[2][0] [5]), .CK(n_59_10), 
      .Q(\buffer[4][2][0] [5]), .QN());
   DFF_X1 \buffer_reg[4][2][0][4]  (.D(\input_filter[2][0] [4]), .CK(n_59_10), 
      .Q(\buffer[4][2][0] [4]), .QN());
   DFF_X1 \buffer_reg[4][2][0][3]  (.D(\input_filter[2][0] [3]), .CK(n_59_10), 
      .Q(\buffer[4][2][0] [3]), .QN());
   DFF_X1 \buffer_reg[4][2][0][2]  (.D(\input_filter[2][0] [2]), .CK(n_59_10), 
      .Q(\buffer[4][2][0] [2]), .QN());
   DFF_X1 \buffer_reg[4][2][0][1]  (.D(\input_filter[2][0] [1]), .CK(n_59_10), 
      .Q(\buffer[4][2][0] [1]), .QN());
   DFF_X1 \buffer_reg[4][2][0][0]  (.D(\input_filter[2][0] [0]), .CK(n_59_10), 
      .Q(\buffer[4][2][0] [0]), .QN());
   DFF_X1 \buffer_reg[5][2][0][15]  (.D(\input_filter[2][0] [15]), .CK(n_59_11), 
      .Q(\buffer[5][2][0] [15]), .QN());
   DFF_X1 \buffer_reg[5][2][0][14]  (.D(\input_filter[2][0] [14]), .CK(n_59_11), 
      .Q(\buffer[5][2][0] [14]), .QN());
   DFF_X1 \buffer_reg[5][2][0][13]  (.D(\input_filter[2][0] [13]), .CK(n_59_11), 
      .Q(\buffer[5][2][0] [13]), .QN());
   DFF_X1 \buffer_reg[5][2][0][12]  (.D(\input_filter[2][0] [12]), .CK(n_59_11), 
      .Q(\buffer[5][2][0] [12]), .QN());
   DFF_X1 \buffer_reg[5][2][0][11]  (.D(\input_filter[2][0] [11]), .CK(n_59_11), 
      .Q(\buffer[5][2][0] [11]), .QN());
   DFF_X1 \buffer_reg[5][2][0][10]  (.D(\input_filter[2][0] [10]), .CK(n_59_11), 
      .Q(\buffer[5][2][0] [10]), .QN());
   DFF_X1 \buffer_reg[5][2][0][9]  (.D(\input_filter[2][0] [9]), .CK(n_59_11), 
      .Q(\buffer[5][2][0] [9]), .QN());
   DFF_X1 \buffer_reg[5][2][0][8]  (.D(\input_filter[2][0] [8]), .CK(n_59_11), 
      .Q(\buffer[5][2][0] [8]), .QN());
   DFF_X1 \buffer_reg[5][2][0][7]  (.D(\input_filter[2][0] [7]), .CK(n_59_11), 
      .Q(\buffer[5][2][0] [7]), .QN());
   DFF_X1 \buffer_reg[5][2][0][6]  (.D(\input_filter[2][0] [6]), .CK(n_59_11), 
      .Q(\buffer[5][2][0] [6]), .QN());
   DFF_X1 \buffer_reg[5][2][0][5]  (.D(\input_filter[2][0] [5]), .CK(n_59_11), 
      .Q(\buffer[5][2][0] [5]), .QN());
   DFF_X1 \buffer_reg[5][2][0][4]  (.D(\input_filter[2][0] [4]), .CK(n_59_11), 
      .Q(\buffer[5][2][0] [4]), .QN());
   DFF_X1 \buffer_reg[5][2][0][3]  (.D(\input_filter[2][0] [3]), .CK(n_59_11), 
      .Q(\buffer[5][2][0] [3]), .QN());
   DFF_X1 \buffer_reg[5][2][0][2]  (.D(\input_filter[2][0] [2]), .CK(n_59_11), 
      .Q(\buffer[5][2][0] [2]), .QN());
   DFF_X1 \buffer_reg[5][2][0][1]  (.D(\input_filter[2][0] [1]), .CK(n_59_11), 
      .Q(\buffer[5][2][0] [1]), .QN());
   DFF_X1 \buffer_reg[5][2][0][0]  (.D(\input_filter[2][0] [0]), .CK(n_59_11), 
      .Q(\buffer[5][2][0] [0]), .QN());
   DFF_X1 \buffer_reg[6][2][0][15]  (.D(\input_filter[2][0] [15]), .CK(n_59_12), 
      .Q(\buffer[6][2][0] [15]), .QN());
   DFF_X1 \buffer_reg[6][2][0][14]  (.D(\input_filter[2][0] [14]), .CK(n_59_12), 
      .Q(\buffer[6][2][0] [14]), .QN());
   DFF_X1 \buffer_reg[6][2][0][13]  (.D(\input_filter[2][0] [13]), .CK(n_59_12), 
      .Q(\buffer[6][2][0] [13]), .QN());
   DFF_X1 \buffer_reg[6][2][0][12]  (.D(\input_filter[2][0] [12]), .CK(n_59_12), 
      .Q(\buffer[6][2][0] [12]), .QN());
   DFF_X1 \buffer_reg[6][2][0][11]  (.D(\input_filter[2][0] [11]), .CK(n_59_12), 
      .Q(\buffer[6][2][0] [11]), .QN());
   DFF_X1 \buffer_reg[6][2][0][10]  (.D(\input_filter[2][0] [10]), .CK(n_59_12), 
      .Q(\buffer[6][2][0] [10]), .QN());
   DFF_X1 \buffer_reg[6][2][0][9]  (.D(\input_filter[2][0] [9]), .CK(n_59_12), 
      .Q(\buffer[6][2][0] [9]), .QN());
   DFF_X1 \buffer_reg[6][2][0][8]  (.D(\input_filter[2][0] [8]), .CK(n_59_12), 
      .Q(\buffer[6][2][0] [8]), .QN());
   DFF_X1 \buffer_reg[6][2][0][7]  (.D(\input_filter[2][0] [7]), .CK(n_59_12), 
      .Q(\buffer[6][2][0] [7]), .QN());
   DFF_X1 \buffer_reg[6][2][0][6]  (.D(\input_filter[2][0] [6]), .CK(n_59_12), 
      .Q(\buffer[6][2][0] [6]), .QN());
   DFF_X1 \buffer_reg[6][2][0][5]  (.D(\input_filter[2][0] [5]), .CK(n_59_12), 
      .Q(\buffer[6][2][0] [5]), .QN());
   DFF_X1 \buffer_reg[6][2][0][4]  (.D(\input_filter[2][0] [4]), .CK(n_59_12), 
      .Q(\buffer[6][2][0] [4]), .QN());
   DFF_X1 \buffer_reg[6][2][0][3]  (.D(\input_filter[2][0] [3]), .CK(n_59_12), 
      .Q(\buffer[6][2][0] [3]), .QN());
   DFF_X1 \buffer_reg[6][2][0][2]  (.D(\input_filter[2][0] [2]), .CK(n_59_12), 
      .Q(\buffer[6][2][0] [2]), .QN());
   DFF_X1 \buffer_reg[6][2][0][1]  (.D(\input_filter[2][0] [1]), .CK(n_59_12), 
      .Q(\buffer[6][2][0] [1]), .QN());
   DFF_X1 \buffer_reg[6][2][0][0]  (.D(\input_filter[2][0] [0]), .CK(n_59_12), 
      .Q(\buffer[6][2][0] [0]), .QN());
   DFF_X1 \buffer_reg[7][2][0][15]  (.D(\input_filter[2][0] [15]), .CK(n_59_13), 
      .Q(\buffer[7][2][0] [15]), .QN());
   DFF_X1 \buffer_reg[7][2][0][14]  (.D(\input_filter[2][0] [14]), .CK(n_59_13), 
      .Q(\buffer[7][2][0] [14]), .QN());
   DFF_X1 \buffer_reg[7][2][0][13]  (.D(\input_filter[2][0] [13]), .CK(n_59_13), 
      .Q(\buffer[7][2][0] [13]), .QN());
   DFF_X1 \buffer_reg[7][2][0][12]  (.D(\input_filter[2][0] [12]), .CK(n_59_13), 
      .Q(\buffer[7][2][0] [12]), .QN());
   DFF_X1 \buffer_reg[7][2][0][11]  (.D(\input_filter[2][0] [11]), .CK(n_59_13), 
      .Q(\buffer[7][2][0] [11]), .QN());
   DFF_X1 \buffer_reg[7][2][0][10]  (.D(\input_filter[2][0] [10]), .CK(n_59_13), 
      .Q(\buffer[7][2][0] [10]), .QN());
   DFF_X1 \buffer_reg[7][2][0][9]  (.D(\input_filter[2][0] [9]), .CK(n_59_13), 
      .Q(\buffer[7][2][0] [9]), .QN());
   DFF_X1 \buffer_reg[7][2][0][8]  (.D(\input_filter[2][0] [8]), .CK(n_59_13), 
      .Q(\buffer[7][2][0] [8]), .QN());
   DFF_X1 \buffer_reg[7][2][0][7]  (.D(\input_filter[2][0] [7]), .CK(n_59_13), 
      .Q(\buffer[7][2][0] [7]), .QN());
   DFF_X1 \buffer_reg[7][2][0][6]  (.D(\input_filter[2][0] [6]), .CK(n_59_13), 
      .Q(\buffer[7][2][0] [6]), .QN());
   DFF_X1 \buffer_reg[7][2][0][5]  (.D(\input_filter[2][0] [5]), .CK(n_59_13), 
      .Q(\buffer[7][2][0] [5]), .QN());
   DFF_X1 \buffer_reg[7][2][0][4]  (.D(\input_filter[2][0] [4]), .CK(n_59_13), 
      .Q(\buffer[7][2][0] [4]), .QN());
   DFF_X1 \buffer_reg[7][2][0][3]  (.D(\input_filter[2][0] [3]), .CK(n_59_13), 
      .Q(\buffer[7][2][0] [3]), .QN());
   DFF_X1 \buffer_reg[7][2][0][2]  (.D(\input_filter[2][0] [2]), .CK(n_59_13), 
      .Q(\buffer[7][2][0] [2]), .QN());
   DFF_X1 \buffer_reg[7][2][0][1]  (.D(\input_filter[2][0] [1]), .CK(n_59_13), 
      .Q(\buffer[7][2][0] [1]), .QN());
   DFF_X1 \buffer_reg[7][2][0][0]  (.D(\input_filter[2][0] [0]), .CK(n_59_13), 
      .Q(\buffer[7][2][0] [0]), .QN());
   DFF_X1 \buffer_reg[8][2][0][15]  (.D(\input_filter[2][0] [15]), .CK(n_59_14), 
      .Q(\buffer[8][2][0] [15]), .QN());
   DFF_X1 \buffer_reg[8][2][0][14]  (.D(\input_filter[2][0] [14]), .CK(n_59_14), 
      .Q(\buffer[8][2][0] [14]), .QN());
   DFF_X1 \buffer_reg[8][2][0][13]  (.D(\input_filter[2][0] [13]), .CK(n_59_14), 
      .Q(\buffer[8][2][0] [13]), .QN());
   DFF_X1 \buffer_reg[8][2][0][12]  (.D(\input_filter[2][0] [12]), .CK(n_59_14), 
      .Q(\buffer[8][2][0] [12]), .QN());
   DFF_X1 \buffer_reg[8][2][0][11]  (.D(\input_filter[2][0] [11]), .CK(n_59_14), 
      .Q(\buffer[8][2][0] [11]), .QN());
   DFF_X1 \buffer_reg[8][2][0][10]  (.D(\input_filter[2][0] [10]), .CK(n_59_14), 
      .Q(\buffer[8][2][0] [10]), .QN());
   DFF_X1 \buffer_reg[8][2][0][9]  (.D(\input_filter[2][0] [9]), .CK(n_59_14), 
      .Q(\buffer[8][2][0] [9]), .QN());
   DFF_X1 \buffer_reg[8][2][0][8]  (.D(\input_filter[2][0] [8]), .CK(n_59_14), 
      .Q(\buffer[8][2][0] [8]), .QN());
   DFF_X1 \buffer_reg[8][2][0][7]  (.D(\input_filter[2][0] [7]), .CK(n_59_14), 
      .Q(\buffer[8][2][0] [7]), .QN());
   DFF_X1 \buffer_reg[8][2][0][6]  (.D(\input_filter[2][0] [6]), .CK(n_59_14), 
      .Q(\buffer[8][2][0] [6]), .QN());
   DFF_X1 \buffer_reg[8][2][0][5]  (.D(\input_filter[2][0] [5]), .CK(n_59_14), 
      .Q(\buffer[8][2][0] [5]), .QN());
   DFF_X1 \buffer_reg[8][2][0][4]  (.D(\input_filter[2][0] [4]), .CK(n_59_14), 
      .Q(\buffer[8][2][0] [4]), .QN());
   DFF_X1 \buffer_reg[8][2][0][3]  (.D(\input_filter[2][0] [3]), .CK(n_59_14), 
      .Q(\buffer[8][2][0] [3]), .QN());
   DFF_X1 \buffer_reg[8][2][0][2]  (.D(\input_filter[2][0] [2]), .CK(n_59_14), 
      .Q(\buffer[8][2][0] [2]), .QN());
   DFF_X1 \buffer_reg[8][2][0][1]  (.D(\input_filter[2][0] [1]), .CK(n_59_14), 
      .Q(\buffer[8][2][0] [1]), .QN());
   DFF_X1 \buffer_reg[8][2][0][0]  (.D(\input_filter[2][0] [0]), .CK(n_59_14), 
      .Q(\buffer[8][2][0] [0]), .QN());
   DFF_X1 \buffer_reg[9][2][0][15]  (.D(\input_filter[2][0] [15]), .CK(n_59_15), 
      .Q(\buffer[9][2][0] [15]), .QN());
   DFF_X1 \buffer_reg[9][2][0][14]  (.D(\input_filter[2][0] [14]), .CK(n_59_15), 
      .Q(\buffer[9][2][0] [14]), .QN());
   DFF_X1 \buffer_reg[9][2][0][13]  (.D(\input_filter[2][0] [13]), .CK(n_59_15), 
      .Q(\buffer[9][2][0] [13]), .QN());
   DFF_X1 \buffer_reg[9][2][0][12]  (.D(\input_filter[2][0] [12]), .CK(n_59_15), 
      .Q(\buffer[9][2][0] [12]), .QN());
   DFF_X1 \buffer_reg[9][2][0][11]  (.D(\input_filter[2][0] [11]), .CK(n_59_15), 
      .Q(\buffer[9][2][0] [11]), .QN());
   DFF_X1 \buffer_reg[9][2][0][10]  (.D(\input_filter[2][0] [10]), .CK(n_59_15), 
      .Q(\buffer[9][2][0] [10]), .QN());
   DFF_X1 \buffer_reg[9][2][0][9]  (.D(\input_filter[2][0] [9]), .CK(n_59_15), 
      .Q(\buffer[9][2][0] [9]), .QN());
   DFF_X1 \buffer_reg[9][2][0][8]  (.D(\input_filter[2][0] [8]), .CK(n_59_15), 
      .Q(\buffer[9][2][0] [8]), .QN());
   DFF_X1 \buffer_reg[9][2][0][7]  (.D(\input_filter[2][0] [7]), .CK(n_59_15), 
      .Q(\buffer[9][2][0] [7]), .QN());
   DFF_X1 \buffer_reg[9][2][0][6]  (.D(\input_filter[2][0] [6]), .CK(n_59_15), 
      .Q(\buffer[9][2][0] [6]), .QN());
   DFF_X1 \buffer_reg[9][2][0][5]  (.D(\input_filter[2][0] [5]), .CK(n_59_15), 
      .Q(\buffer[9][2][0] [5]), .QN());
   DFF_X1 \buffer_reg[9][2][0][4]  (.D(\input_filter[2][0] [4]), .CK(n_59_15), 
      .Q(\buffer[9][2][0] [4]), .QN());
   DFF_X1 \buffer_reg[9][2][0][3]  (.D(\input_filter[2][0] [3]), .CK(n_59_15), 
      .Q(\buffer[9][2][0] [3]), .QN());
   DFF_X1 \buffer_reg[9][2][0][2]  (.D(\input_filter[2][0] [2]), .CK(n_59_15), 
      .Q(\buffer[9][2][0] [2]), .QN());
   DFF_X1 \buffer_reg[9][2][0][1]  (.D(\input_filter[2][0] [1]), .CK(n_59_15), 
      .Q(\buffer[9][2][0] [1]), .QN());
   DFF_X1 \buffer_reg[9][2][0][0]  (.D(\input_filter[2][0] [0]), .CK(n_59_15), 
      .Q(\buffer[9][2][0] [0]), .QN());
   DFF_X1 \buffer_reg[10][2][0][15]  (.D(\input_filter[2][0] [15]), .CK(n_59_6), 
      .Q(\buffer[10][2][0] [15]), .QN());
   DFF_X1 \buffer_reg[10][2][0][14]  (.D(\input_filter[2][0] [14]), .CK(n_59_6), 
      .Q(\buffer[10][2][0] [14]), .QN());
   DFF_X1 \buffer_reg[10][2][0][13]  (.D(\input_filter[2][0] [13]), .CK(n_59_6), 
      .Q(\buffer[10][2][0] [13]), .QN());
   DFF_X1 \buffer_reg[10][2][0][12]  (.D(\input_filter[2][0] [12]), .CK(n_59_6), 
      .Q(\buffer[10][2][0] [12]), .QN());
   DFF_X1 \buffer_reg[10][2][0][11]  (.D(\input_filter[2][0] [11]), .CK(n_59_6), 
      .Q(\buffer[10][2][0] [11]), .QN());
   DFF_X1 \buffer_reg[10][2][0][10]  (.D(\input_filter[2][0] [10]), .CK(n_59_6), 
      .Q(\buffer[10][2][0] [10]), .QN());
   DFF_X1 \buffer_reg[10][2][0][9]  (.D(\input_filter[2][0] [9]), .CK(n_59_6), 
      .Q(\buffer[10][2][0] [9]), .QN());
   DFF_X1 \buffer_reg[10][2][0][8]  (.D(\input_filter[2][0] [8]), .CK(n_59_6), 
      .Q(\buffer[10][2][0] [8]), .QN());
   DFF_X1 \buffer_reg[10][2][0][7]  (.D(\input_filter[2][0] [7]), .CK(n_59_6), 
      .Q(\buffer[10][2][0] [7]), .QN());
   DFF_X1 \buffer_reg[10][2][0][6]  (.D(\input_filter[2][0] [6]), .CK(n_59_6), 
      .Q(\buffer[10][2][0] [6]), .QN());
   DFF_X1 \buffer_reg[10][2][0][5]  (.D(\input_filter[2][0] [5]), .CK(n_59_6), 
      .Q(\buffer[10][2][0] [5]), .QN());
   DFF_X1 \buffer_reg[10][2][0][4]  (.D(\input_filter[2][0] [4]), .CK(n_59_6), 
      .Q(\buffer[10][2][0] [4]), .QN());
   DFF_X1 \buffer_reg[10][2][0][3]  (.D(\input_filter[2][0] [3]), .CK(n_59_6), 
      .Q(\buffer[10][2][0] [3]), .QN());
   DFF_X1 \buffer_reg[10][2][0][2]  (.D(\input_filter[2][0] [2]), .CK(n_59_6), 
      .Q(\buffer[10][2][0] [2]), .QN());
   DFF_X1 \buffer_reg[10][2][0][1]  (.D(\input_filter[2][0] [1]), .CK(n_59_6), 
      .Q(\buffer[10][2][0] [1]), .QN());
   DFF_X1 \buffer_reg[10][2][0][0]  (.D(\input_filter[2][0] [0]), .CK(n_59_6), 
      .Q(\buffer[10][2][0] [0]), .QN());
   DFF_X1 \buffer_reg[11][2][0][15]  (.D(\input_filter[2][0] [15]), .CK(n_59_1), 
      .Q(\buffer[11][2][0] [15]), .QN());
   DFF_X1 \buffer_reg[11][2][0][14]  (.D(\input_filter[2][0] [14]), .CK(n_59_1), 
      .Q(\buffer[11][2][0] [14]), .QN());
   DFF_X1 \buffer_reg[11][2][0][13]  (.D(\input_filter[2][0] [13]), .CK(n_59_1), 
      .Q(\buffer[11][2][0] [13]), .QN());
   DFF_X1 \buffer_reg[11][2][0][12]  (.D(\input_filter[2][0] [12]), .CK(n_59_1), 
      .Q(\buffer[11][2][0] [12]), .QN());
   DFF_X1 \buffer_reg[11][2][0][11]  (.D(\input_filter[2][0] [11]), .CK(n_59_1), 
      .Q(\buffer[11][2][0] [11]), .QN());
   DFF_X1 \buffer_reg[11][2][0][10]  (.D(\input_filter[2][0] [10]), .CK(n_59_1), 
      .Q(\buffer[11][2][0] [10]), .QN());
   DFF_X1 \buffer_reg[11][2][0][9]  (.D(\input_filter[2][0] [9]), .CK(n_59_1), 
      .Q(\buffer[11][2][0] [9]), .QN());
   DFF_X1 \buffer_reg[11][2][0][8]  (.D(\input_filter[2][0] [8]), .CK(n_59_1), 
      .Q(\buffer[11][2][0] [8]), .QN());
   DFF_X1 \buffer_reg[11][2][0][7]  (.D(\input_filter[2][0] [7]), .CK(n_59_1), 
      .Q(\buffer[11][2][0] [7]), .QN());
   DFF_X1 \buffer_reg[11][2][0][6]  (.D(\input_filter[2][0] [6]), .CK(n_59_1), 
      .Q(\buffer[11][2][0] [6]), .QN());
   DFF_X1 \buffer_reg[11][2][0][5]  (.D(\input_filter[2][0] [5]), .CK(n_59_1), 
      .Q(\buffer[11][2][0] [5]), .QN());
   DFF_X1 \buffer_reg[11][2][0][4]  (.D(\input_filter[2][0] [4]), .CK(n_59_1), 
      .Q(\buffer[11][2][0] [4]), .QN());
   DFF_X1 \buffer_reg[11][2][0][3]  (.D(\input_filter[2][0] [3]), .CK(n_59_1), 
      .Q(\buffer[11][2][0] [3]), .QN());
   DFF_X1 \buffer_reg[11][2][0][2]  (.D(\input_filter[2][0] [2]), .CK(n_59_1), 
      .Q(\buffer[11][2][0] [2]), .QN());
   DFF_X1 \buffer_reg[11][2][0][1]  (.D(\input_filter[2][0] [1]), .CK(n_59_1), 
      .Q(\buffer[11][2][0] [1]), .QN());
   DFF_X1 \buffer_reg[11][2][0][0]  (.D(\input_filter[2][0] [0]), .CK(n_59_1), 
      .Q(\buffer[11][2][0] [0]), .QN());
   DFF_X1 \buffer_reg[12][2][0][15]  (.D(\input_filter[2][0] [15]), .CK(n_59_2), 
      .Q(\buffer[12][2][0] [15]), .QN());
   DFF_X1 \buffer_reg[12][2][0][14]  (.D(\input_filter[2][0] [14]), .CK(n_59_2), 
      .Q(\buffer[12][2][0] [14]), .QN());
   DFF_X1 \buffer_reg[12][2][0][13]  (.D(\input_filter[2][0] [13]), .CK(n_59_2), 
      .Q(\buffer[12][2][0] [13]), .QN());
   DFF_X1 \buffer_reg[12][2][0][12]  (.D(\input_filter[2][0] [12]), .CK(n_59_2), 
      .Q(\buffer[12][2][0] [12]), .QN());
   DFF_X1 \buffer_reg[12][2][0][11]  (.D(\input_filter[2][0] [11]), .CK(n_59_2), 
      .Q(\buffer[12][2][0] [11]), .QN());
   DFF_X1 \buffer_reg[12][2][0][10]  (.D(\input_filter[2][0] [10]), .CK(n_59_2), 
      .Q(\buffer[12][2][0] [10]), .QN());
   DFF_X1 \buffer_reg[12][2][0][9]  (.D(\input_filter[2][0] [9]), .CK(n_59_2), 
      .Q(\buffer[12][2][0] [9]), .QN());
   DFF_X1 \buffer_reg[12][2][0][8]  (.D(\input_filter[2][0] [8]), .CK(n_59_2), 
      .Q(\buffer[12][2][0] [8]), .QN());
   DFF_X1 \buffer_reg[12][2][0][7]  (.D(\input_filter[2][0] [7]), .CK(n_59_2), 
      .Q(\buffer[12][2][0] [7]), .QN());
   DFF_X1 \buffer_reg[12][2][0][6]  (.D(\input_filter[2][0] [6]), .CK(n_59_2), 
      .Q(\buffer[12][2][0] [6]), .QN());
   DFF_X1 \buffer_reg[12][2][0][5]  (.D(\input_filter[2][0] [5]), .CK(n_59_2), 
      .Q(\buffer[12][2][0] [5]), .QN());
   DFF_X1 \buffer_reg[12][2][0][4]  (.D(\input_filter[2][0] [4]), .CK(n_59_2), 
      .Q(\buffer[12][2][0] [4]), .QN());
   DFF_X1 \buffer_reg[12][2][0][3]  (.D(\input_filter[2][0] [3]), .CK(n_59_2), 
      .Q(\buffer[12][2][0] [3]), .QN());
   DFF_X1 \buffer_reg[12][2][0][2]  (.D(\input_filter[2][0] [2]), .CK(n_59_2), 
      .Q(\buffer[12][2][0] [2]), .QN());
   DFF_X1 \buffer_reg[12][2][0][1]  (.D(\input_filter[2][0] [1]), .CK(n_59_2), 
      .Q(\buffer[12][2][0] [1]), .QN());
   DFF_X1 \buffer_reg[12][2][0][0]  (.D(\input_filter[2][0] [0]), .CK(n_59_2), 
      .Q(\buffer[12][2][0] [0]), .QN());
   DFF_X1 \buffer_reg[13][2][0][15]  (.D(\input_filter[2][0] [15]), .CK(n_59_3), 
      .Q(\buffer[13][2][0] [15]), .QN());
   DFF_X1 \buffer_reg[13][2][0][14]  (.D(\input_filter[2][0] [14]), .CK(n_59_3), 
      .Q(\buffer[13][2][0] [14]), .QN());
   DFF_X1 \buffer_reg[13][2][0][13]  (.D(\input_filter[2][0] [13]), .CK(n_59_3), 
      .Q(\buffer[13][2][0] [13]), .QN());
   DFF_X1 \buffer_reg[13][2][0][12]  (.D(\input_filter[2][0] [12]), .CK(n_59_3), 
      .Q(\buffer[13][2][0] [12]), .QN());
   DFF_X1 \buffer_reg[13][2][0][11]  (.D(\input_filter[2][0] [11]), .CK(n_59_3), 
      .Q(\buffer[13][2][0] [11]), .QN());
   DFF_X1 \buffer_reg[13][2][0][10]  (.D(\input_filter[2][0] [10]), .CK(n_59_3), 
      .Q(\buffer[13][2][0] [10]), .QN());
   DFF_X1 \buffer_reg[13][2][0][9]  (.D(\input_filter[2][0] [9]), .CK(n_59_3), 
      .Q(\buffer[13][2][0] [9]), .QN());
   DFF_X1 \buffer_reg[13][2][0][8]  (.D(\input_filter[2][0] [8]), .CK(n_59_3), 
      .Q(\buffer[13][2][0] [8]), .QN());
   DFF_X1 \buffer_reg[13][2][0][7]  (.D(\input_filter[2][0] [7]), .CK(n_59_3), 
      .Q(\buffer[13][2][0] [7]), .QN());
   DFF_X1 \buffer_reg[13][2][0][6]  (.D(\input_filter[2][0] [6]), .CK(n_59_3), 
      .Q(\buffer[13][2][0] [6]), .QN());
   DFF_X1 \buffer_reg[13][2][0][5]  (.D(\input_filter[2][0] [5]), .CK(n_59_3), 
      .Q(\buffer[13][2][0] [5]), .QN());
   DFF_X1 \buffer_reg[13][2][0][4]  (.D(\input_filter[2][0] [4]), .CK(n_59_3), 
      .Q(\buffer[13][2][0] [4]), .QN());
   DFF_X1 \buffer_reg[13][2][0][3]  (.D(\input_filter[2][0] [3]), .CK(n_59_3), 
      .Q(\buffer[13][2][0] [3]), .QN());
   DFF_X1 \buffer_reg[13][2][0][2]  (.D(\input_filter[2][0] [2]), .CK(n_59_3), 
      .Q(\buffer[13][2][0] [2]), .QN());
   DFF_X1 \buffer_reg[13][2][0][1]  (.D(\input_filter[2][0] [1]), .CK(n_59_3), 
      .Q(\buffer[13][2][0] [1]), .QN());
   DFF_X1 \buffer_reg[13][2][0][0]  (.D(\input_filter[2][0] [0]), .CK(n_59_3), 
      .Q(\buffer[13][2][0] [0]), .QN());
   DFF_X1 \buffer_reg[14][2][0][15]  (.D(\input_filter[2][0] [15]), .CK(n_59_4), 
      .Q(\buffer[14][2][0] [15]), .QN());
   DFF_X1 \buffer_reg[14][2][0][14]  (.D(\input_filter[2][0] [14]), .CK(n_59_4), 
      .Q(\buffer[14][2][0] [14]), .QN());
   DFF_X1 \buffer_reg[14][2][0][13]  (.D(\input_filter[2][0] [13]), .CK(n_59_4), 
      .Q(\buffer[14][2][0] [13]), .QN());
   DFF_X1 \buffer_reg[14][2][0][12]  (.D(\input_filter[2][0] [12]), .CK(n_59_4), 
      .Q(\buffer[14][2][0] [12]), .QN());
   DFF_X1 \buffer_reg[14][2][0][11]  (.D(\input_filter[2][0] [11]), .CK(n_59_4), 
      .Q(\buffer[14][2][0] [11]), .QN());
   DFF_X1 \buffer_reg[14][2][0][10]  (.D(\input_filter[2][0] [10]), .CK(n_59_4), 
      .Q(\buffer[14][2][0] [10]), .QN());
   DFF_X1 \buffer_reg[14][2][0][9]  (.D(\input_filter[2][0] [9]), .CK(n_59_4), 
      .Q(\buffer[14][2][0] [9]), .QN());
   DFF_X1 \buffer_reg[14][2][0][8]  (.D(\input_filter[2][0] [8]), .CK(n_59_4), 
      .Q(\buffer[14][2][0] [8]), .QN());
   DFF_X1 \buffer_reg[14][2][0][7]  (.D(\input_filter[2][0] [7]), .CK(n_59_4), 
      .Q(\buffer[14][2][0] [7]), .QN());
   DFF_X1 \buffer_reg[14][2][0][6]  (.D(\input_filter[2][0] [6]), .CK(n_59_4), 
      .Q(\buffer[14][2][0] [6]), .QN());
   DFF_X1 \buffer_reg[14][2][0][5]  (.D(\input_filter[2][0] [5]), .CK(n_59_4), 
      .Q(\buffer[14][2][0] [5]), .QN());
   DFF_X1 \buffer_reg[14][2][0][4]  (.D(\input_filter[2][0] [4]), .CK(n_59_4), 
      .Q(\buffer[14][2][0] [4]), .QN());
   DFF_X1 \buffer_reg[14][2][0][3]  (.D(\input_filter[2][0] [3]), .CK(n_59_4), 
      .Q(\buffer[14][2][0] [3]), .QN());
   DFF_X1 \buffer_reg[14][2][0][2]  (.D(\input_filter[2][0] [2]), .CK(n_59_4), 
      .Q(\buffer[14][2][0] [2]), .QN());
   DFF_X1 \buffer_reg[14][2][0][1]  (.D(\input_filter[2][0] [1]), .CK(n_59_4), 
      .Q(\buffer[14][2][0] [1]), .QN());
   DFF_X1 \buffer_reg[14][2][0][0]  (.D(\input_filter[2][0] [0]), .CK(n_59_4), 
      .Q(\buffer[14][2][0] [0]), .QN());
   DFF_X1 \buffer_reg[15][2][0][15]  (.D(\input_filter[2][0] [15]), .CK(n_59_5), 
      .Q(\buffer[15][2][0] [15]), .QN());
   DFF_X1 \buffer_reg[15][2][0][14]  (.D(\input_filter[2][0] [14]), .CK(n_59_5), 
      .Q(\buffer[15][2][0] [14]), .QN());
   DFF_X1 \buffer_reg[15][2][0][13]  (.D(\input_filter[2][0] [13]), .CK(n_59_5), 
      .Q(\buffer[15][2][0] [13]), .QN());
   DFF_X1 \buffer_reg[15][2][0][12]  (.D(\input_filter[2][0] [12]), .CK(n_59_5), 
      .Q(\buffer[15][2][0] [12]), .QN());
   DFF_X1 \buffer_reg[15][2][0][11]  (.D(\input_filter[2][0] [11]), .CK(n_59_5), 
      .Q(\buffer[15][2][0] [11]), .QN());
   DFF_X1 \buffer_reg[15][2][0][10]  (.D(\input_filter[2][0] [10]), .CK(n_59_5), 
      .Q(\buffer[15][2][0] [10]), .QN());
   DFF_X1 \buffer_reg[15][2][0][9]  (.D(\input_filter[2][0] [9]), .CK(n_59_5), 
      .Q(\buffer[15][2][0] [9]), .QN());
   DFF_X1 \buffer_reg[15][2][0][8]  (.D(\input_filter[2][0] [8]), .CK(n_59_5), 
      .Q(\buffer[15][2][0] [8]), .QN());
   DFF_X1 \buffer_reg[15][2][0][7]  (.D(\input_filter[2][0] [7]), .CK(n_59_5), 
      .Q(\buffer[15][2][0] [7]), .QN());
   DFF_X1 \buffer_reg[15][2][0][6]  (.D(\input_filter[2][0] [6]), .CK(n_59_5), 
      .Q(\buffer[15][2][0] [6]), .QN());
   DFF_X1 \buffer_reg[15][2][0][5]  (.D(\input_filter[2][0] [5]), .CK(n_59_5), 
      .Q(\buffer[15][2][0] [5]), .QN());
   DFF_X1 \buffer_reg[15][2][0][4]  (.D(\input_filter[2][0] [4]), .CK(n_59_5), 
      .Q(\buffer[15][2][0] [4]), .QN());
   DFF_X1 \buffer_reg[15][2][0][3]  (.D(\input_filter[2][0] [3]), .CK(n_59_5), 
      .Q(\buffer[15][2][0] [3]), .QN());
   DFF_X1 \buffer_reg[15][2][0][2]  (.D(\input_filter[2][0] [2]), .CK(n_59_5), 
      .Q(\buffer[15][2][0] [2]), .QN());
   DFF_X1 \buffer_reg[15][2][0][1]  (.D(\input_filter[2][0] [1]), .CK(n_59_5), 
      .Q(\buffer[15][2][0] [1]), .QN());
   DFF_X1 \buffer_reg[15][2][0][0]  (.D(\input_filter[2][0] [0]), .CK(n_59_5), 
      .Q(\buffer[15][2][0] [0]), .QN());
   DFF_X1 \buffer_reg[12][2][1][15]  (.D(\input_filter[2][1] [15]), .CK(n_59_2), 
      .Q(\buffer[12][2][1] [15]), .QN());
   DFF_X1 \buffer_reg[12][2][1][14]  (.D(\input_filter[2][1] [14]), .CK(n_59_2), 
      .Q(\buffer[12][2][1] [14]), .QN());
   DFF_X1 \buffer_reg[12][2][1][13]  (.D(\input_filter[2][1] [13]), .CK(n_59_2), 
      .Q(\buffer[12][2][1] [13]), .QN());
   DFF_X1 \buffer_reg[12][2][1][12]  (.D(\input_filter[2][1] [12]), .CK(n_59_2), 
      .Q(\buffer[12][2][1] [12]), .QN());
   DFF_X1 \buffer_reg[12][2][1][11]  (.D(\input_filter[2][1] [11]), .CK(n_59_2), 
      .Q(\buffer[12][2][1] [11]), .QN());
   DFF_X1 \buffer_reg[12][2][1][10]  (.D(\input_filter[2][1] [10]), .CK(n_59_2), 
      .Q(\buffer[12][2][1] [10]), .QN());
   DFF_X1 \buffer_reg[12][2][1][9]  (.D(\input_filter[2][1] [9]), .CK(n_59_2), 
      .Q(\buffer[12][2][1] [9]), .QN());
   DFF_X1 \buffer_reg[12][2][1][8]  (.D(\input_filter[2][1] [8]), .CK(n_59_2), 
      .Q(\buffer[12][2][1] [8]), .QN());
   DFF_X1 \buffer_reg[12][2][1][7]  (.D(\input_filter[2][1] [7]), .CK(n_59_2), 
      .Q(\buffer[12][2][1] [7]), .QN());
   DFF_X1 \buffer_reg[12][2][1][6]  (.D(\input_filter[2][1] [6]), .CK(n_59_2), 
      .Q(\buffer[12][2][1] [6]), .QN());
   DFF_X1 \buffer_reg[12][2][1][5]  (.D(\input_filter[2][1] [5]), .CK(n_59_2), 
      .Q(\buffer[12][2][1] [5]), .QN());
   DFF_X1 \buffer_reg[12][2][1][4]  (.D(\input_filter[2][1] [4]), .CK(n_59_2), 
      .Q(\buffer[12][2][1] [4]), .QN());
   DFF_X1 \buffer_reg[12][2][1][3]  (.D(\input_filter[2][1] [3]), .CK(n_59_2), 
      .Q(\buffer[12][2][1] [3]), .QN());
   DFF_X1 \buffer_reg[12][2][1][2]  (.D(\input_filter[2][1] [2]), .CK(n_59_2), 
      .Q(\buffer[12][2][1] [2]), .QN());
   DFF_X1 \buffer_reg[12][2][1][1]  (.D(\input_filter[2][1] [1]), .CK(n_59_2), 
      .Q(\buffer[12][2][1] [1]), .QN());
   DFF_X1 \buffer_reg[12][2][1][0]  (.D(\input_filter[2][1] [0]), .CK(n_59_2), 
      .Q(\buffer[12][2][1] [0]), .QN());
   DFF_X1 \buffer_reg[0][2][1][15]  (.D(\input_filter[2][1] [15]), .CK(n_59_0), 
      .Q(\buffer[0][2][1] [15]), .QN());
   DFF_X1 \buffer_reg[0][2][1][14]  (.D(\input_filter[2][1] [14]), .CK(n_59_0), 
      .Q(\buffer[0][2][1] [14]), .QN());
   DFF_X1 \buffer_reg[0][2][1][13]  (.D(\input_filter[2][1] [13]), .CK(n_59_0), 
      .Q(\buffer[0][2][1] [13]), .QN());
   DFF_X1 \buffer_reg[0][2][1][12]  (.D(\input_filter[2][1] [12]), .CK(n_59_0), 
      .Q(\buffer[0][2][1] [12]), .QN());
   DFF_X1 \buffer_reg[0][2][1][11]  (.D(\input_filter[2][1] [11]), .CK(n_59_0), 
      .Q(\buffer[0][2][1] [11]), .QN());
   DFF_X1 \buffer_reg[0][2][1][10]  (.D(\input_filter[2][1] [10]), .CK(n_59_0), 
      .Q(\buffer[0][2][1] [10]), .QN());
   DFF_X1 \buffer_reg[0][2][1][9]  (.D(\input_filter[2][1] [9]), .CK(n_59_0), 
      .Q(\buffer[0][2][1] [9]), .QN());
   DFF_X1 \buffer_reg[0][2][1][8]  (.D(\input_filter[2][1] [8]), .CK(n_59_0), 
      .Q(\buffer[0][2][1] [8]), .QN());
   DFF_X1 \buffer_reg[0][2][1][7]  (.D(\input_filter[2][1] [7]), .CK(n_59_0), 
      .Q(\buffer[0][2][1] [7]), .QN());
   DFF_X1 \buffer_reg[0][2][1][6]  (.D(\input_filter[2][1] [6]), .CK(n_59_0), 
      .Q(\buffer[0][2][1] [6]), .QN());
   DFF_X1 \buffer_reg[0][2][1][5]  (.D(\input_filter[2][1] [5]), .CK(n_59_0), 
      .Q(\buffer[0][2][1] [5]), .QN());
   DFF_X1 \buffer_reg[0][2][1][4]  (.D(\input_filter[2][1] [4]), .CK(n_59_0), 
      .Q(\buffer[0][2][1] [4]), .QN());
   DFF_X1 \buffer_reg[0][2][1][3]  (.D(\input_filter[2][1] [3]), .CK(n_59_0), 
      .Q(\buffer[0][2][1] [3]), .QN());
   DFF_X1 \buffer_reg[0][2][1][2]  (.D(\input_filter[2][1] [2]), .CK(n_59_0), 
      .Q(\buffer[0][2][1] [2]), .QN());
   DFF_X1 \buffer_reg[0][2][1][1]  (.D(\input_filter[2][1] [1]), .CK(n_59_0), 
      .Q(\buffer[0][2][1] [1]), .QN());
   DFF_X1 \buffer_reg[0][2][1][0]  (.D(\input_filter[2][1] [0]), .CK(n_59_0), 
      .Q(\buffer[0][2][1] [0]), .QN());
   DFF_X1 \buffer_reg[1][2][1][15]  (.D(\input_filter[2][1] [15]), .CK(n_59_7), 
      .Q(\buffer[1][2][1] [15]), .QN());
   DFF_X1 \buffer_reg[1][2][1][14]  (.D(\input_filter[2][1] [14]), .CK(n_59_7), 
      .Q(\buffer[1][2][1] [14]), .QN());
   DFF_X1 \buffer_reg[1][2][1][13]  (.D(\input_filter[2][1] [13]), .CK(n_59_7), 
      .Q(\buffer[1][2][1] [13]), .QN());
   DFF_X1 \buffer_reg[1][2][1][12]  (.D(\input_filter[2][1] [12]), .CK(n_59_7), 
      .Q(\buffer[1][2][1] [12]), .QN());
   DFF_X1 \buffer_reg[1][2][1][11]  (.D(\input_filter[2][1] [11]), .CK(n_59_7), 
      .Q(\buffer[1][2][1] [11]), .QN());
   DFF_X1 \buffer_reg[1][2][1][10]  (.D(\input_filter[2][1] [10]), .CK(n_59_7), 
      .Q(\buffer[1][2][1] [10]), .QN());
   DFF_X1 \buffer_reg[1][2][1][9]  (.D(\input_filter[2][1] [9]), .CK(n_59_7), 
      .Q(\buffer[1][2][1] [9]), .QN());
   DFF_X1 \buffer_reg[1][2][1][8]  (.D(\input_filter[2][1] [8]), .CK(n_59_7), 
      .Q(\buffer[1][2][1] [8]), .QN());
   DFF_X1 \buffer_reg[1][2][1][7]  (.D(\input_filter[2][1] [7]), .CK(n_59_7), 
      .Q(\buffer[1][2][1] [7]), .QN());
   DFF_X1 \buffer_reg[1][2][1][6]  (.D(\input_filter[2][1] [6]), .CK(n_59_7), 
      .Q(\buffer[1][2][1] [6]), .QN());
   DFF_X1 \buffer_reg[1][2][1][5]  (.D(\input_filter[2][1] [5]), .CK(n_59_7), 
      .Q(\buffer[1][2][1] [5]), .QN());
   DFF_X1 \buffer_reg[1][2][1][4]  (.D(\input_filter[2][1] [4]), .CK(n_59_7), 
      .Q(\buffer[1][2][1] [4]), .QN());
   DFF_X1 \buffer_reg[1][2][1][3]  (.D(\input_filter[2][1] [3]), .CK(n_59_7), 
      .Q(\buffer[1][2][1] [3]), .QN());
   DFF_X1 \buffer_reg[1][2][1][2]  (.D(\input_filter[2][1] [2]), .CK(n_59_7), 
      .Q(\buffer[1][2][1] [2]), .QN());
   DFF_X1 \buffer_reg[1][2][1][1]  (.D(\input_filter[2][1] [1]), .CK(n_59_7), 
      .Q(\buffer[1][2][1] [1]), .QN());
   DFF_X1 \buffer_reg[1][2][1][0]  (.D(\input_filter[2][1] [0]), .CK(n_59_7), 
      .Q(\buffer[1][2][1] [0]), .QN());
   DFF_X1 \buffer_reg[2][2][1][15]  (.D(\input_filter[2][1] [15]), .CK(n_59_8), 
      .Q(\buffer[2][2][1] [15]), .QN());
   DFF_X1 \buffer_reg[2][2][1][14]  (.D(\input_filter[2][1] [14]), .CK(n_59_8), 
      .Q(\buffer[2][2][1] [14]), .QN());
   DFF_X1 \buffer_reg[2][2][1][13]  (.D(\input_filter[2][1] [13]), .CK(n_59_8), 
      .Q(\buffer[2][2][1] [13]), .QN());
   DFF_X1 \buffer_reg[2][2][1][12]  (.D(\input_filter[2][1] [12]), .CK(n_59_8), 
      .Q(\buffer[2][2][1] [12]), .QN());
   DFF_X1 \buffer_reg[2][2][1][11]  (.D(\input_filter[2][1] [11]), .CK(n_59_8), 
      .Q(\buffer[2][2][1] [11]), .QN());
   DFF_X1 \buffer_reg[2][2][1][10]  (.D(\input_filter[2][1] [10]), .CK(n_59_8), 
      .Q(\buffer[2][2][1] [10]), .QN());
   DFF_X1 \buffer_reg[2][2][1][9]  (.D(\input_filter[2][1] [9]), .CK(n_59_8), 
      .Q(\buffer[2][2][1] [9]), .QN());
   DFF_X1 \buffer_reg[2][2][1][8]  (.D(\input_filter[2][1] [8]), .CK(n_59_8), 
      .Q(\buffer[2][2][1] [8]), .QN());
   DFF_X1 \buffer_reg[2][2][1][7]  (.D(\input_filter[2][1] [7]), .CK(n_59_8), 
      .Q(\buffer[2][2][1] [7]), .QN());
   DFF_X1 \buffer_reg[2][2][1][6]  (.D(\input_filter[2][1] [6]), .CK(n_59_8), 
      .Q(\buffer[2][2][1] [6]), .QN());
   DFF_X1 \buffer_reg[2][2][1][5]  (.D(\input_filter[2][1] [5]), .CK(n_59_8), 
      .Q(\buffer[2][2][1] [5]), .QN());
   DFF_X1 \buffer_reg[2][2][1][4]  (.D(\input_filter[2][1] [4]), .CK(n_59_8), 
      .Q(\buffer[2][2][1] [4]), .QN());
   DFF_X1 \buffer_reg[2][2][1][3]  (.D(\input_filter[2][1] [3]), .CK(n_59_8), 
      .Q(\buffer[2][2][1] [3]), .QN());
   DFF_X1 \buffer_reg[2][2][1][2]  (.D(\input_filter[2][1] [2]), .CK(n_59_8), 
      .Q(\buffer[2][2][1] [2]), .QN());
   DFF_X1 \buffer_reg[2][2][1][1]  (.D(\input_filter[2][1] [1]), .CK(n_59_8), 
      .Q(\buffer[2][2][1] [1]), .QN());
   DFF_X1 \buffer_reg[2][2][1][0]  (.D(\input_filter[2][1] [0]), .CK(n_59_8), 
      .Q(\buffer[2][2][1] [0]), .QN());
   DFF_X1 \buffer_reg[3][2][1][15]  (.D(\input_filter[2][1] [15]), .CK(n_59_9), 
      .Q(\buffer[3][2][1] [15]), .QN());
   DFF_X1 \buffer_reg[3][2][1][14]  (.D(\input_filter[2][1] [14]), .CK(n_59_9), 
      .Q(\buffer[3][2][1] [14]), .QN());
   DFF_X1 \buffer_reg[3][2][1][13]  (.D(\input_filter[2][1] [13]), .CK(n_59_9), 
      .Q(\buffer[3][2][1] [13]), .QN());
   DFF_X1 \buffer_reg[3][2][1][12]  (.D(\input_filter[2][1] [12]), .CK(n_59_9), 
      .Q(\buffer[3][2][1] [12]), .QN());
   DFF_X1 \buffer_reg[3][2][1][11]  (.D(\input_filter[2][1] [11]), .CK(n_59_9), 
      .Q(\buffer[3][2][1] [11]), .QN());
   DFF_X1 \buffer_reg[3][2][1][10]  (.D(\input_filter[2][1] [10]), .CK(n_59_9), 
      .Q(\buffer[3][2][1] [10]), .QN());
   DFF_X1 \buffer_reg[3][2][1][9]  (.D(\input_filter[2][1] [9]), .CK(n_59_9), 
      .Q(\buffer[3][2][1] [9]), .QN());
   DFF_X1 \buffer_reg[3][2][1][8]  (.D(\input_filter[2][1] [8]), .CK(n_59_9), 
      .Q(\buffer[3][2][1] [8]), .QN());
   DFF_X1 \buffer_reg[3][2][1][7]  (.D(\input_filter[2][1] [7]), .CK(n_59_9), 
      .Q(\buffer[3][2][1] [7]), .QN());
   DFF_X1 \buffer_reg[3][2][1][6]  (.D(\input_filter[2][1] [6]), .CK(n_59_9), 
      .Q(\buffer[3][2][1] [6]), .QN());
   DFF_X1 \buffer_reg[3][2][1][5]  (.D(\input_filter[2][1] [5]), .CK(n_59_9), 
      .Q(\buffer[3][2][1] [5]), .QN());
   DFF_X1 \buffer_reg[3][2][1][4]  (.D(\input_filter[2][1] [4]), .CK(n_59_9), 
      .Q(\buffer[3][2][1] [4]), .QN());
   DFF_X1 \buffer_reg[3][2][1][3]  (.D(\input_filter[2][1] [3]), .CK(n_59_9), 
      .Q(\buffer[3][2][1] [3]), .QN());
   DFF_X1 \buffer_reg[3][2][1][2]  (.D(\input_filter[2][1] [2]), .CK(n_59_9), 
      .Q(\buffer[3][2][1] [2]), .QN());
   DFF_X1 \buffer_reg[3][2][1][1]  (.D(\input_filter[2][1] [1]), .CK(n_59_9), 
      .Q(\buffer[3][2][1] [1]), .QN());
   DFF_X1 \buffer_reg[3][2][1][0]  (.D(\input_filter[2][1] [0]), .CK(n_59_9), 
      .Q(\buffer[3][2][1] [0]), .QN());
   DFF_X1 \buffer_reg[4][2][1][15]  (.D(\input_filter[2][1] [15]), .CK(n_59_10), 
      .Q(\buffer[4][2][1] [15]), .QN());
   DFF_X1 \buffer_reg[4][2][1][14]  (.D(\input_filter[2][1] [14]), .CK(n_59_10), 
      .Q(\buffer[4][2][1] [14]), .QN());
   DFF_X1 \buffer_reg[4][2][1][13]  (.D(\input_filter[2][1] [13]), .CK(n_59_10), 
      .Q(\buffer[4][2][1] [13]), .QN());
   DFF_X1 \buffer_reg[4][2][1][12]  (.D(\input_filter[2][1] [12]), .CK(n_59_10), 
      .Q(\buffer[4][2][1] [12]), .QN());
   DFF_X1 \buffer_reg[4][2][1][11]  (.D(\input_filter[2][1] [11]), .CK(n_59_10), 
      .Q(\buffer[4][2][1] [11]), .QN());
   DFF_X1 \buffer_reg[4][2][1][10]  (.D(\input_filter[2][1] [10]), .CK(n_59_10), 
      .Q(\buffer[4][2][1] [10]), .QN());
   DFF_X1 \buffer_reg[4][2][1][9]  (.D(\input_filter[2][1] [9]), .CK(n_59_10), 
      .Q(\buffer[4][2][1] [9]), .QN());
   DFF_X1 \buffer_reg[4][2][1][8]  (.D(\input_filter[2][1] [8]), .CK(n_59_10), 
      .Q(\buffer[4][2][1] [8]), .QN());
   DFF_X1 \buffer_reg[4][2][1][7]  (.D(\input_filter[2][1] [7]), .CK(n_59_10), 
      .Q(\buffer[4][2][1] [7]), .QN());
   DFF_X1 \buffer_reg[4][2][1][6]  (.D(\input_filter[2][1] [6]), .CK(n_59_10), 
      .Q(\buffer[4][2][1] [6]), .QN());
   DFF_X1 \buffer_reg[4][2][1][5]  (.D(\input_filter[2][1] [5]), .CK(n_59_10), 
      .Q(\buffer[4][2][1] [5]), .QN());
   DFF_X1 \buffer_reg[4][2][1][4]  (.D(\input_filter[2][1] [4]), .CK(n_59_10), 
      .Q(\buffer[4][2][1] [4]), .QN());
   DFF_X1 \buffer_reg[4][2][1][3]  (.D(\input_filter[2][1] [3]), .CK(n_59_10), 
      .Q(\buffer[4][2][1] [3]), .QN());
   DFF_X1 \buffer_reg[4][2][1][2]  (.D(\input_filter[2][1] [2]), .CK(n_59_10), 
      .Q(\buffer[4][2][1] [2]), .QN());
   DFF_X1 \buffer_reg[4][2][1][1]  (.D(\input_filter[2][1] [1]), .CK(n_59_10), 
      .Q(\buffer[4][2][1] [1]), .QN());
   DFF_X1 \buffer_reg[4][2][1][0]  (.D(\input_filter[2][1] [0]), .CK(n_59_10), 
      .Q(\buffer[4][2][1] [0]), .QN());
   DFF_X1 \buffer_reg[5][2][1][15]  (.D(\input_filter[2][1] [15]), .CK(n_59_11), 
      .Q(\buffer[5][2][1] [15]), .QN());
   DFF_X1 \buffer_reg[5][2][1][14]  (.D(\input_filter[2][1] [14]), .CK(n_59_11), 
      .Q(\buffer[5][2][1] [14]), .QN());
   DFF_X1 \buffer_reg[5][2][1][13]  (.D(\input_filter[2][1] [13]), .CK(n_59_11), 
      .Q(\buffer[5][2][1] [13]), .QN());
   DFF_X1 \buffer_reg[5][2][1][12]  (.D(\input_filter[2][1] [12]), .CK(n_59_11), 
      .Q(\buffer[5][2][1] [12]), .QN());
   DFF_X1 \buffer_reg[5][2][1][11]  (.D(\input_filter[2][1] [11]), .CK(n_59_11), 
      .Q(\buffer[5][2][1] [11]), .QN());
   DFF_X1 \buffer_reg[5][2][1][10]  (.D(\input_filter[2][1] [10]), .CK(n_59_11), 
      .Q(\buffer[5][2][1] [10]), .QN());
   DFF_X1 \buffer_reg[5][2][1][9]  (.D(\input_filter[2][1] [9]), .CK(n_59_11), 
      .Q(\buffer[5][2][1] [9]), .QN());
   DFF_X1 \buffer_reg[5][2][1][8]  (.D(\input_filter[2][1] [8]), .CK(n_59_11), 
      .Q(\buffer[5][2][1] [8]), .QN());
   DFF_X1 \buffer_reg[5][2][1][7]  (.D(\input_filter[2][1] [7]), .CK(n_59_11), 
      .Q(\buffer[5][2][1] [7]), .QN());
   DFF_X1 \buffer_reg[5][2][1][6]  (.D(\input_filter[2][1] [6]), .CK(n_59_11), 
      .Q(\buffer[5][2][1] [6]), .QN());
   DFF_X1 \buffer_reg[5][2][1][5]  (.D(\input_filter[2][1] [5]), .CK(n_59_11), 
      .Q(\buffer[5][2][1] [5]), .QN());
   DFF_X1 \buffer_reg[5][2][1][4]  (.D(\input_filter[2][1] [4]), .CK(n_59_11), 
      .Q(\buffer[5][2][1] [4]), .QN());
   DFF_X1 \buffer_reg[5][2][1][3]  (.D(\input_filter[2][1] [3]), .CK(n_59_11), 
      .Q(\buffer[5][2][1] [3]), .QN());
   DFF_X1 \buffer_reg[5][2][1][2]  (.D(\input_filter[2][1] [2]), .CK(n_59_11), 
      .Q(\buffer[5][2][1] [2]), .QN());
   DFF_X1 \buffer_reg[5][2][1][1]  (.D(\input_filter[2][1] [1]), .CK(n_59_11), 
      .Q(\buffer[5][2][1] [1]), .QN());
   DFF_X1 \buffer_reg[5][2][1][0]  (.D(\input_filter[2][1] [0]), .CK(n_59_11), 
      .Q(\buffer[5][2][1] [0]), .QN());
   DFF_X1 \buffer_reg[6][2][1][15]  (.D(\input_filter[2][1] [15]), .CK(n_59_12), 
      .Q(\buffer[6][2][1] [15]), .QN());
   DFF_X1 \buffer_reg[6][2][1][14]  (.D(\input_filter[2][1] [14]), .CK(n_59_12), 
      .Q(\buffer[6][2][1] [14]), .QN());
   DFF_X1 \buffer_reg[6][2][1][13]  (.D(\input_filter[2][1] [13]), .CK(n_59_12), 
      .Q(\buffer[6][2][1] [13]), .QN());
   DFF_X1 \buffer_reg[6][2][1][12]  (.D(\input_filter[2][1] [12]), .CK(n_59_12), 
      .Q(\buffer[6][2][1] [12]), .QN());
   DFF_X1 \buffer_reg[6][2][1][11]  (.D(\input_filter[2][1] [11]), .CK(n_59_12), 
      .Q(\buffer[6][2][1] [11]), .QN());
   DFF_X1 \buffer_reg[6][2][1][10]  (.D(\input_filter[2][1] [10]), .CK(n_59_12), 
      .Q(\buffer[6][2][1] [10]), .QN());
   DFF_X1 \buffer_reg[6][2][1][9]  (.D(\input_filter[2][1] [9]), .CK(n_59_12), 
      .Q(\buffer[6][2][1] [9]), .QN());
   DFF_X1 \buffer_reg[6][2][1][8]  (.D(\input_filter[2][1] [8]), .CK(n_59_12), 
      .Q(\buffer[6][2][1] [8]), .QN());
   DFF_X1 \buffer_reg[6][2][1][7]  (.D(\input_filter[2][1] [7]), .CK(n_59_12), 
      .Q(\buffer[6][2][1] [7]), .QN());
   DFF_X1 \buffer_reg[6][2][1][6]  (.D(\input_filter[2][1] [6]), .CK(n_59_12), 
      .Q(\buffer[6][2][1] [6]), .QN());
   DFF_X1 \buffer_reg[6][2][1][5]  (.D(\input_filter[2][1] [5]), .CK(n_59_12), 
      .Q(\buffer[6][2][1] [5]), .QN());
   DFF_X1 \buffer_reg[6][2][1][4]  (.D(\input_filter[2][1] [4]), .CK(n_59_12), 
      .Q(\buffer[6][2][1] [4]), .QN());
   DFF_X1 \buffer_reg[6][2][1][3]  (.D(\input_filter[2][1] [3]), .CK(n_59_12), 
      .Q(\buffer[6][2][1] [3]), .QN());
   DFF_X1 \buffer_reg[6][2][1][2]  (.D(\input_filter[2][1] [2]), .CK(n_59_12), 
      .Q(\buffer[6][2][1] [2]), .QN());
   DFF_X1 \buffer_reg[6][2][1][1]  (.D(\input_filter[2][1] [1]), .CK(n_59_12), 
      .Q(\buffer[6][2][1] [1]), .QN());
   DFF_X1 \buffer_reg[6][2][1][0]  (.D(\input_filter[2][1] [0]), .CK(n_59_12), 
      .Q(\buffer[6][2][1] [0]), .QN());
   DFF_X1 \buffer_reg[7][2][1][15]  (.D(\input_filter[2][1] [15]), .CK(n_59_13), 
      .Q(\buffer[7][2][1] [15]), .QN());
   DFF_X1 \buffer_reg[7][2][1][14]  (.D(\input_filter[2][1] [14]), .CK(n_59_13), 
      .Q(\buffer[7][2][1] [14]), .QN());
   DFF_X1 \buffer_reg[7][2][1][13]  (.D(\input_filter[2][1] [13]), .CK(n_59_13), 
      .Q(\buffer[7][2][1] [13]), .QN());
   DFF_X1 \buffer_reg[7][2][1][12]  (.D(\input_filter[2][1] [12]), .CK(n_59_13), 
      .Q(\buffer[7][2][1] [12]), .QN());
   DFF_X1 \buffer_reg[7][2][1][11]  (.D(\input_filter[2][1] [11]), .CK(n_59_13), 
      .Q(\buffer[7][2][1] [11]), .QN());
   DFF_X1 \buffer_reg[7][2][1][10]  (.D(\input_filter[2][1] [10]), .CK(n_59_13), 
      .Q(\buffer[7][2][1] [10]), .QN());
   DFF_X1 \buffer_reg[7][2][1][9]  (.D(\input_filter[2][1] [9]), .CK(n_59_13), 
      .Q(\buffer[7][2][1] [9]), .QN());
   DFF_X1 \buffer_reg[7][2][1][8]  (.D(\input_filter[2][1] [8]), .CK(n_59_13), 
      .Q(\buffer[7][2][1] [8]), .QN());
   DFF_X1 \buffer_reg[7][2][1][7]  (.D(\input_filter[2][1] [7]), .CK(n_59_13), 
      .Q(\buffer[7][2][1] [7]), .QN());
   DFF_X1 \buffer_reg[7][2][1][6]  (.D(\input_filter[2][1] [6]), .CK(n_59_13), 
      .Q(\buffer[7][2][1] [6]), .QN());
   DFF_X1 \buffer_reg[7][2][1][5]  (.D(\input_filter[2][1] [5]), .CK(n_59_13), 
      .Q(\buffer[7][2][1] [5]), .QN());
   DFF_X1 \buffer_reg[7][2][1][4]  (.D(\input_filter[2][1] [4]), .CK(n_59_13), 
      .Q(\buffer[7][2][1] [4]), .QN());
   DFF_X1 \buffer_reg[7][2][1][3]  (.D(\input_filter[2][1] [3]), .CK(n_59_13), 
      .Q(\buffer[7][2][1] [3]), .QN());
   DFF_X1 \buffer_reg[7][2][1][2]  (.D(\input_filter[2][1] [2]), .CK(n_59_13), 
      .Q(\buffer[7][2][1] [2]), .QN());
   DFF_X1 \buffer_reg[7][2][1][1]  (.D(\input_filter[2][1] [1]), .CK(n_59_13), 
      .Q(\buffer[7][2][1] [1]), .QN());
   DFF_X1 \buffer_reg[7][2][1][0]  (.D(\input_filter[2][1] [0]), .CK(n_59_13), 
      .Q(\buffer[7][2][1] [0]), .QN());
   DFF_X1 \buffer_reg[8][2][1][15]  (.D(\input_filter[2][1] [15]), .CK(n_59_14), 
      .Q(\buffer[8][2][1] [15]), .QN());
   DFF_X1 \buffer_reg[8][2][1][14]  (.D(\input_filter[2][1] [14]), .CK(n_59_14), 
      .Q(\buffer[8][2][1] [14]), .QN());
   DFF_X1 \buffer_reg[8][2][1][13]  (.D(\input_filter[2][1] [13]), .CK(n_59_14), 
      .Q(\buffer[8][2][1] [13]), .QN());
   DFF_X1 \buffer_reg[8][2][1][12]  (.D(\input_filter[2][1] [12]), .CK(n_59_14), 
      .Q(\buffer[8][2][1] [12]), .QN());
   DFF_X1 \buffer_reg[8][2][1][11]  (.D(\input_filter[2][1] [11]), .CK(n_59_14), 
      .Q(\buffer[8][2][1] [11]), .QN());
   DFF_X1 \buffer_reg[8][2][1][10]  (.D(\input_filter[2][1] [10]), .CK(n_59_14), 
      .Q(\buffer[8][2][1] [10]), .QN());
   DFF_X1 \buffer_reg[8][2][1][9]  (.D(\input_filter[2][1] [9]), .CK(n_59_14), 
      .Q(\buffer[8][2][1] [9]), .QN());
   DFF_X1 \buffer_reg[8][2][1][8]  (.D(\input_filter[2][1] [8]), .CK(n_59_14), 
      .Q(\buffer[8][2][1] [8]), .QN());
   DFF_X1 \buffer_reg[8][2][1][7]  (.D(\input_filter[2][1] [7]), .CK(n_59_14), 
      .Q(\buffer[8][2][1] [7]), .QN());
   DFF_X1 \buffer_reg[8][2][1][6]  (.D(\input_filter[2][1] [6]), .CK(n_59_14), 
      .Q(\buffer[8][2][1] [6]), .QN());
   DFF_X1 \buffer_reg[8][2][1][5]  (.D(\input_filter[2][1] [5]), .CK(n_59_14), 
      .Q(\buffer[8][2][1] [5]), .QN());
   DFF_X1 \buffer_reg[8][2][1][4]  (.D(\input_filter[2][1] [4]), .CK(n_59_14), 
      .Q(\buffer[8][2][1] [4]), .QN());
   DFF_X1 \buffer_reg[8][2][1][3]  (.D(\input_filter[2][1] [3]), .CK(n_59_14), 
      .Q(\buffer[8][2][1] [3]), .QN());
   DFF_X1 \buffer_reg[8][2][1][2]  (.D(\input_filter[2][1] [2]), .CK(n_59_14), 
      .Q(\buffer[8][2][1] [2]), .QN());
   DFF_X1 \buffer_reg[8][2][1][1]  (.D(\input_filter[2][1] [1]), .CK(n_59_14), 
      .Q(\buffer[8][2][1] [1]), .QN());
   DFF_X1 \buffer_reg[8][2][1][0]  (.D(\input_filter[2][1] [0]), .CK(n_59_14), 
      .Q(\buffer[8][2][1] [0]), .QN());
   DFF_X1 \buffer_reg[9][2][1][15]  (.D(\input_filter[2][1] [15]), .CK(n_59_15), 
      .Q(\buffer[9][2][1] [15]), .QN());
   DFF_X1 \buffer_reg[9][2][1][14]  (.D(\input_filter[2][1] [14]), .CK(n_59_15), 
      .Q(\buffer[9][2][1] [14]), .QN());
   DFF_X1 \buffer_reg[9][2][1][13]  (.D(\input_filter[2][1] [13]), .CK(n_59_15), 
      .Q(\buffer[9][2][1] [13]), .QN());
   DFF_X1 \buffer_reg[9][2][1][12]  (.D(\input_filter[2][1] [12]), .CK(n_59_15), 
      .Q(\buffer[9][2][1] [12]), .QN());
   DFF_X1 \buffer_reg[9][2][1][11]  (.D(\input_filter[2][1] [11]), .CK(n_59_15), 
      .Q(\buffer[9][2][1] [11]), .QN());
   DFF_X1 \buffer_reg[9][2][1][10]  (.D(\input_filter[2][1] [10]), .CK(n_59_15), 
      .Q(\buffer[9][2][1] [10]), .QN());
   DFF_X1 \buffer_reg[9][2][1][9]  (.D(\input_filter[2][1] [9]), .CK(n_59_15), 
      .Q(\buffer[9][2][1] [9]), .QN());
   DFF_X1 \buffer_reg[9][2][1][8]  (.D(\input_filter[2][1] [8]), .CK(n_59_15), 
      .Q(\buffer[9][2][1] [8]), .QN());
   DFF_X1 \buffer_reg[9][2][1][7]  (.D(\input_filter[2][1] [7]), .CK(n_59_15), 
      .Q(\buffer[9][2][1] [7]), .QN());
   DFF_X1 \buffer_reg[9][2][1][6]  (.D(\input_filter[2][1] [6]), .CK(n_59_15), 
      .Q(\buffer[9][2][1] [6]), .QN());
   DFF_X1 \buffer_reg[9][2][1][5]  (.D(\input_filter[2][1] [5]), .CK(n_59_15), 
      .Q(\buffer[9][2][1] [5]), .QN());
   DFF_X1 \buffer_reg[9][2][1][4]  (.D(\input_filter[2][1] [4]), .CK(n_59_15), 
      .Q(\buffer[9][2][1] [4]), .QN());
   DFF_X1 \buffer_reg[9][2][1][3]  (.D(\input_filter[2][1] [3]), .CK(n_59_15), 
      .Q(\buffer[9][2][1] [3]), .QN());
   DFF_X1 \buffer_reg[9][2][1][2]  (.D(\input_filter[2][1] [2]), .CK(n_59_15), 
      .Q(\buffer[9][2][1] [2]), .QN());
   DFF_X1 \buffer_reg[9][2][1][1]  (.D(\input_filter[2][1] [1]), .CK(n_59_15), 
      .Q(\buffer[9][2][1] [1]), .QN());
   DFF_X1 \buffer_reg[9][2][1][0]  (.D(\input_filter[2][1] [0]), .CK(n_59_15), 
      .Q(\buffer[9][2][1] [0]), .QN());
   DFF_X1 \buffer_reg[10][2][1][15]  (.D(\input_filter[2][1] [15]), .CK(n_59_6), 
      .Q(\buffer[10][2][1] [15]), .QN());
   DFF_X1 \buffer_reg[10][2][1][14]  (.D(\input_filter[2][1] [14]), .CK(n_59_6), 
      .Q(\buffer[10][2][1] [14]), .QN());
   DFF_X1 \buffer_reg[10][2][1][13]  (.D(\input_filter[2][1] [13]), .CK(n_59_6), 
      .Q(\buffer[10][2][1] [13]), .QN());
   DFF_X1 \buffer_reg[10][2][1][12]  (.D(\input_filter[2][1] [12]), .CK(n_59_6), 
      .Q(\buffer[10][2][1] [12]), .QN());
   DFF_X1 \buffer_reg[10][2][1][11]  (.D(\input_filter[2][1] [11]), .CK(n_59_6), 
      .Q(\buffer[10][2][1] [11]), .QN());
   DFF_X1 \buffer_reg[10][2][1][10]  (.D(\input_filter[2][1] [10]), .CK(n_59_6), 
      .Q(\buffer[10][2][1] [10]), .QN());
   DFF_X1 \buffer_reg[10][2][1][9]  (.D(\input_filter[2][1] [9]), .CK(n_59_6), 
      .Q(\buffer[10][2][1] [9]), .QN());
   DFF_X1 \buffer_reg[10][2][1][8]  (.D(\input_filter[2][1] [8]), .CK(n_59_6), 
      .Q(\buffer[10][2][1] [8]), .QN());
   DFF_X1 \buffer_reg[10][2][1][7]  (.D(\input_filter[2][1] [7]), .CK(n_59_6), 
      .Q(\buffer[10][2][1] [7]), .QN());
   DFF_X1 \buffer_reg[10][2][1][6]  (.D(\input_filter[2][1] [6]), .CK(n_59_6), 
      .Q(\buffer[10][2][1] [6]), .QN());
   DFF_X1 \buffer_reg[10][2][1][5]  (.D(\input_filter[2][1] [5]), .CK(n_59_6), 
      .Q(\buffer[10][2][1] [5]), .QN());
   DFF_X1 \buffer_reg[10][2][1][4]  (.D(\input_filter[2][1] [4]), .CK(n_59_6), 
      .Q(\buffer[10][2][1] [4]), .QN());
   DFF_X1 \buffer_reg[10][2][1][3]  (.D(\input_filter[2][1] [3]), .CK(n_59_6), 
      .Q(\buffer[10][2][1] [3]), .QN());
   DFF_X1 \buffer_reg[10][2][1][2]  (.D(\input_filter[2][1] [2]), .CK(n_59_6), 
      .Q(\buffer[10][2][1] [2]), .QN());
   DFF_X1 \buffer_reg[10][2][1][1]  (.D(\input_filter[2][1] [1]), .CK(n_59_6), 
      .Q(\buffer[10][2][1] [1]), .QN());
   DFF_X1 \buffer_reg[10][2][1][0]  (.D(\input_filter[2][1] [0]), .CK(n_59_6), 
      .Q(\buffer[10][2][1] [0]), .QN());
   DFF_X1 \buffer_reg[11][2][1][15]  (.D(\input_filter[2][1] [15]), .CK(n_59_1), 
      .Q(\buffer[11][2][1] [15]), .QN());
   DFF_X1 \buffer_reg[11][2][1][14]  (.D(\input_filter[2][1] [14]), .CK(n_59_1), 
      .Q(\buffer[11][2][1] [14]), .QN());
   DFF_X1 \buffer_reg[11][2][1][13]  (.D(\input_filter[2][1] [13]), .CK(n_59_1), 
      .Q(\buffer[11][2][1] [13]), .QN());
   DFF_X1 \buffer_reg[11][2][1][12]  (.D(\input_filter[2][1] [12]), .CK(n_59_1), 
      .Q(\buffer[11][2][1] [12]), .QN());
   DFF_X1 \buffer_reg[11][2][1][11]  (.D(\input_filter[2][1] [11]), .CK(n_59_1), 
      .Q(\buffer[11][2][1] [11]), .QN());
   DFF_X1 \buffer_reg[11][2][1][10]  (.D(\input_filter[2][1] [10]), .CK(n_59_1), 
      .Q(\buffer[11][2][1] [10]), .QN());
   DFF_X1 \buffer_reg[11][2][1][9]  (.D(\input_filter[2][1] [9]), .CK(n_59_1), 
      .Q(\buffer[11][2][1] [9]), .QN());
   DFF_X1 \buffer_reg[11][2][1][8]  (.D(\input_filter[2][1] [8]), .CK(n_59_1), 
      .Q(\buffer[11][2][1] [8]), .QN());
   DFF_X1 \buffer_reg[11][2][1][7]  (.D(\input_filter[2][1] [7]), .CK(n_59_1), 
      .Q(\buffer[11][2][1] [7]), .QN());
   DFF_X1 \buffer_reg[11][2][1][6]  (.D(\input_filter[2][1] [6]), .CK(n_59_1), 
      .Q(\buffer[11][2][1] [6]), .QN());
   DFF_X1 \buffer_reg[11][2][1][5]  (.D(\input_filter[2][1] [5]), .CK(n_59_1), 
      .Q(\buffer[11][2][1] [5]), .QN());
   DFF_X1 \buffer_reg[11][2][1][4]  (.D(\input_filter[2][1] [4]), .CK(n_59_1), 
      .Q(\buffer[11][2][1] [4]), .QN());
   DFF_X1 \buffer_reg[11][2][1][3]  (.D(\input_filter[2][1] [3]), .CK(n_59_1), 
      .Q(\buffer[11][2][1] [3]), .QN());
   DFF_X1 \buffer_reg[11][2][1][2]  (.D(\input_filter[2][1] [2]), .CK(n_59_1), 
      .Q(\buffer[11][2][1] [2]), .QN());
   DFF_X1 \buffer_reg[11][2][1][1]  (.D(\input_filter[2][1] [1]), .CK(n_59_1), 
      .Q(\buffer[11][2][1] [1]), .QN());
   DFF_X1 \buffer_reg[11][2][1][0]  (.D(\input_filter[2][1] [0]), .CK(n_59_1), 
      .Q(\buffer[11][2][1] [0]), .QN());
   DFF_X1 \buffer_reg[13][2][1][15]  (.D(\input_filter[2][1] [15]), .CK(n_59_3), 
      .Q(\buffer[13][2][1] [15]), .QN());
   DFF_X1 \buffer_reg[13][2][1][14]  (.D(\input_filter[2][1] [14]), .CK(n_59_3), 
      .Q(\buffer[13][2][1] [14]), .QN());
   DFF_X1 \buffer_reg[13][2][1][13]  (.D(\input_filter[2][1] [13]), .CK(n_59_3), 
      .Q(\buffer[13][2][1] [13]), .QN());
   DFF_X1 \buffer_reg[13][2][1][12]  (.D(\input_filter[2][1] [12]), .CK(n_59_3), 
      .Q(\buffer[13][2][1] [12]), .QN());
   DFF_X1 \buffer_reg[13][2][1][11]  (.D(\input_filter[2][1] [11]), .CK(n_59_3), 
      .Q(\buffer[13][2][1] [11]), .QN());
   DFF_X1 \buffer_reg[13][2][1][10]  (.D(\input_filter[2][1] [10]), .CK(n_59_3), 
      .Q(\buffer[13][2][1] [10]), .QN());
   DFF_X1 \buffer_reg[13][2][1][9]  (.D(\input_filter[2][1] [9]), .CK(n_59_3), 
      .Q(\buffer[13][2][1] [9]), .QN());
   DFF_X1 \buffer_reg[13][2][1][8]  (.D(\input_filter[2][1] [8]), .CK(n_59_3), 
      .Q(\buffer[13][2][1] [8]), .QN());
   DFF_X1 \buffer_reg[13][2][1][7]  (.D(\input_filter[2][1] [7]), .CK(n_59_3), 
      .Q(\buffer[13][2][1] [7]), .QN());
   DFF_X1 \buffer_reg[13][2][1][6]  (.D(\input_filter[2][1] [6]), .CK(n_59_3), 
      .Q(\buffer[13][2][1] [6]), .QN());
   DFF_X1 \buffer_reg[13][2][1][5]  (.D(\input_filter[2][1] [5]), .CK(n_59_3), 
      .Q(\buffer[13][2][1] [5]), .QN());
   DFF_X1 \buffer_reg[13][2][1][4]  (.D(\input_filter[2][1] [4]), .CK(n_59_3), 
      .Q(\buffer[13][2][1] [4]), .QN());
   DFF_X1 \buffer_reg[13][2][1][3]  (.D(\input_filter[2][1] [3]), .CK(n_59_3), 
      .Q(\buffer[13][2][1] [3]), .QN());
   DFF_X1 \buffer_reg[13][2][1][2]  (.D(\input_filter[2][1] [2]), .CK(n_59_3), 
      .Q(\buffer[13][2][1] [2]), .QN());
   DFF_X1 \buffer_reg[13][2][1][1]  (.D(\input_filter[2][1] [1]), .CK(n_59_3), 
      .Q(\buffer[13][2][1] [1]), .QN());
   DFF_X1 \buffer_reg[13][2][1][0]  (.D(\input_filter[2][1] [0]), .CK(n_59_3), 
      .Q(\buffer[13][2][1] [0]), .QN());
   DFF_X1 \buffer_reg[14][2][1][15]  (.D(\input_filter[2][1] [15]), .CK(n_59_4), 
      .Q(\buffer[14][2][1] [15]), .QN());
   DFF_X1 \buffer_reg[14][2][1][14]  (.D(\input_filter[2][1] [14]), .CK(n_59_4), 
      .Q(\buffer[14][2][1] [14]), .QN());
   DFF_X1 \buffer_reg[14][2][1][13]  (.D(\input_filter[2][1] [13]), .CK(n_59_4), 
      .Q(\buffer[14][2][1] [13]), .QN());
   DFF_X1 \buffer_reg[14][2][1][12]  (.D(\input_filter[2][1] [12]), .CK(n_59_4), 
      .Q(\buffer[14][2][1] [12]), .QN());
   DFF_X1 \buffer_reg[14][2][1][11]  (.D(\input_filter[2][1] [11]), .CK(n_59_4), 
      .Q(\buffer[14][2][1] [11]), .QN());
   DFF_X1 \buffer_reg[14][2][1][10]  (.D(\input_filter[2][1] [10]), .CK(n_59_4), 
      .Q(\buffer[14][2][1] [10]), .QN());
   DFF_X1 \buffer_reg[14][2][1][9]  (.D(\input_filter[2][1] [9]), .CK(n_59_4), 
      .Q(\buffer[14][2][1] [9]), .QN());
   DFF_X1 \buffer_reg[14][2][1][8]  (.D(\input_filter[2][1] [8]), .CK(n_59_4), 
      .Q(\buffer[14][2][1] [8]), .QN());
   DFF_X1 \buffer_reg[14][2][1][7]  (.D(\input_filter[2][1] [7]), .CK(n_59_4), 
      .Q(\buffer[14][2][1] [7]), .QN());
   DFF_X1 \buffer_reg[14][2][1][6]  (.D(\input_filter[2][1] [6]), .CK(n_59_4), 
      .Q(\buffer[14][2][1] [6]), .QN());
   DFF_X1 \buffer_reg[14][2][1][5]  (.D(\input_filter[2][1] [5]), .CK(n_59_4), 
      .Q(\buffer[14][2][1] [5]), .QN());
   DFF_X1 \buffer_reg[14][2][1][4]  (.D(\input_filter[2][1] [4]), .CK(n_59_4), 
      .Q(\buffer[14][2][1] [4]), .QN());
   DFF_X1 \buffer_reg[14][2][1][3]  (.D(\input_filter[2][1] [3]), .CK(n_59_4), 
      .Q(\buffer[14][2][1] [3]), .QN());
   DFF_X1 \buffer_reg[14][2][1][2]  (.D(\input_filter[2][1] [2]), .CK(n_59_4), 
      .Q(\buffer[14][2][1] [2]), .QN());
   DFF_X1 \buffer_reg[14][2][1][1]  (.D(\input_filter[2][1] [1]), .CK(n_59_4), 
      .Q(\buffer[14][2][1] [1]), .QN());
   DFF_X1 \buffer_reg[14][2][1][0]  (.D(\input_filter[2][1] [0]), .CK(n_59_4), 
      .Q(\buffer[14][2][1] [0]), .QN());
   DFF_X1 \buffer_reg[15][2][1][15]  (.D(\input_filter[2][1] [15]), .CK(n_59_5), 
      .Q(\buffer[15][2][1] [15]), .QN());
   DFF_X1 \buffer_reg[15][2][1][14]  (.D(\input_filter[2][1] [14]), .CK(n_59_5), 
      .Q(\buffer[15][2][1] [14]), .QN());
   DFF_X1 \buffer_reg[15][2][1][13]  (.D(\input_filter[2][1] [13]), .CK(n_59_5), 
      .Q(\buffer[15][2][1] [13]), .QN());
   DFF_X1 \buffer_reg[15][2][1][12]  (.D(\input_filter[2][1] [12]), .CK(n_59_5), 
      .Q(\buffer[15][2][1] [12]), .QN());
   DFF_X1 \buffer_reg[15][2][1][11]  (.D(\input_filter[2][1] [11]), .CK(n_59_5), 
      .Q(\buffer[15][2][1] [11]), .QN());
   DFF_X1 \buffer_reg[15][2][1][10]  (.D(\input_filter[2][1] [10]), .CK(n_59_5), 
      .Q(\buffer[15][2][1] [10]), .QN());
   DFF_X1 \buffer_reg[15][2][1][9]  (.D(\input_filter[2][1] [9]), .CK(n_59_5), 
      .Q(\buffer[15][2][1] [9]), .QN());
   DFF_X1 \buffer_reg[15][2][1][8]  (.D(\input_filter[2][1] [8]), .CK(n_59_5), 
      .Q(\buffer[15][2][1] [8]), .QN());
   DFF_X1 \buffer_reg[15][2][1][7]  (.D(\input_filter[2][1] [7]), .CK(n_59_5), 
      .Q(\buffer[15][2][1] [7]), .QN());
   DFF_X1 \buffer_reg[15][2][1][6]  (.D(\input_filter[2][1] [6]), .CK(n_59_5), 
      .Q(\buffer[15][2][1] [6]), .QN());
   DFF_X1 \buffer_reg[15][2][1][5]  (.D(\input_filter[2][1] [5]), .CK(n_59_5), 
      .Q(\buffer[15][2][1] [5]), .QN());
   DFF_X1 \buffer_reg[15][2][1][4]  (.D(\input_filter[2][1] [4]), .CK(n_59_5), 
      .Q(\buffer[15][2][1] [4]), .QN());
   DFF_X1 \buffer_reg[15][2][1][3]  (.D(\input_filter[2][1] [3]), .CK(n_59_5), 
      .Q(\buffer[15][2][1] [3]), .QN());
   DFF_X1 \buffer_reg[15][2][1][2]  (.D(\input_filter[2][1] [2]), .CK(n_59_5), 
      .Q(\buffer[15][2][1] [2]), .QN());
   DFF_X1 \buffer_reg[15][2][1][1]  (.D(\input_filter[2][1] [1]), .CK(n_59_5), 
      .Q(\buffer[15][2][1] [1]), .QN());
   DFF_X1 \buffer_reg[15][2][1][0]  (.D(\input_filter[2][1] [0]), .CK(n_59_5), 
      .Q(\buffer[15][2][1] [0]), .QN());
   CLKGATETST_X1 \clk_gate_buffer_reg[0][1][4]_reg  (.CK(read), .E(n_0), 
      .SE(1'b0), .GCK(n_59_0));
   CLKGATETST_X1 \clk_gate_buffer_reg[11][1][4]_reg  (.CK(read), .E(n_11), 
      .SE(1'b0), .GCK(n_59_1));
   CLKGATETST_X1 \clk_gate_buffer_reg[12][1][4]_reg  (.CK(read), .E(n_12), 
      .SE(1'b0), .GCK(n_59_2));
   CLKGATETST_X1 \clk_gate_buffer_reg[13][1][4]_reg  (.CK(read), .E(n_13), 
      .SE(1'b0), .GCK(n_59_3));
   CLKGATETST_X1 \clk_gate_buffer_reg[14][1][4]_reg  (.CK(read), .E(n_14), 
      .SE(1'b0), .GCK(n_59_4));
   CLKGATETST_X1 \clk_gate_buffer_reg[15][1][4]_reg  (.CK(read), .E(n_15), 
      .SE(1'b0), .GCK(n_59_5));
   CLKGATETST_X1 \clk_gate_buffer_reg[1][2][0]_reg  (.CK(read), .E(n_1), 
      .SE(1'b0), .GCK(n_59_7));
   CLKGATETST_X1 \clk_gate_buffer_reg[2][2][0]_reg  (.CK(read), .E(n_2), 
      .SE(1'b0), .GCK(n_59_8));
   CLKGATETST_X1 \clk_gate_buffer_reg[3][2][0]_reg  (.CK(read), .E(n_3), 
      .SE(1'b0), .GCK(n_59_9));
   CLKGATETST_X1 \clk_gate_buffer_reg[4][2][0]_reg  (.CK(read), .E(n_4), 
      .SE(1'b0), .GCK(n_59_10));
   CLKGATETST_X1 \clk_gate_buffer_reg[5][2][0]_reg  (.CK(read), .E(n_5), 
      .SE(1'b0), .GCK(n_59_11));
   CLKGATETST_X1 \clk_gate_buffer_reg[6][2][0]_reg  (.CK(read), .E(n_6), 
      .SE(1'b0), .GCK(n_59_12));
   CLKGATETST_X1 \clk_gate_buffer_reg[7][2][0]_reg  (.CK(read), .E(n_7), 
      .SE(1'b0), .GCK(n_59_13));
   CLKGATETST_X1 \clk_gate_buffer_reg[8][2][0]_reg  (.CK(read), .E(n_8), 
      .SE(1'b0), .GCK(n_59_14));
   CLKGATETST_X1 \clk_gate_buffer_reg[9][2][0]_reg  (.CK(read), .E(n_9), 
      .SE(1'b0), .GCK(n_59_15));
   CLKGATETST_X1 \clk_gate_buffer_reg[10][2][0]_reg  (.CK(read), .E(n_10), 
      .SE(1'b0), .GCK(n_59_6));
   NOR3_X1 i_1_0_0 (.A1(n_1_0_0), .A2(index_buffer[1]), .A3(index_buffer[2]), 
      .ZN(n_0));
   NOR3_X1 i_1_0_1 (.A1(n_1_0_1), .A2(index_buffer[1]), .A3(index_buffer[2]), 
      .ZN(n_1));
   NOR2_X1 i_1_0_2 (.A1(n_1_0_2), .A2(n_1_0_0), .ZN(n_2));
   NOR2_X1 i_1_0_3 (.A1(n_1_0_2), .A2(n_1_0_1), .ZN(n_3));
   NOR2_X1 i_1_0_4 (.A1(n_1_0_3), .A2(n_1_0_0), .ZN(n_4));
   NOR2_X1 i_1_0_5 (.A1(n_1_0_3), .A2(n_1_0_1), .ZN(n_5));
   NOR2_X1 i_1_0_6 (.A1(n_1_0_5), .A2(n_1_0_0), .ZN(n_6));
   NAND3_X1 i_1_0_7 (.A1(n_1_0_7), .A2(n_1_0_11), .A3(n_1_0_13), .ZN(n_1_0_0));
   NOR2_X1 i_1_0_8 (.A1(n_1_0_5), .A2(n_1_0_1), .ZN(n_7));
   NAND3_X1 i_1_0_9 (.A1(n_1_0_7), .A2(n_1_0_13), .A3(index_buffer[0]), .ZN(
      n_1_0_1));
   NOR3_X1 i_1_0_10 (.A1(n_1_0_4), .A2(index_buffer[1]), .A3(index_buffer[2]), 
      .ZN(n_8));
   NOR3_X1 i_1_0_11 (.A1(n_1_0_6), .A2(index_buffer[1]), .A3(index_buffer[2]), 
      .ZN(n_9));
   NOR2_X1 i_1_0_12 (.A1(n_1_0_4), .A2(n_1_0_2), .ZN(n_10));
   NOR2_X1 i_1_0_13 (.A1(n_1_0_6), .A2(n_1_0_2), .ZN(n_11));
   OR2_X1 i_1_0_14 (.A1(n_1_0_12), .A2(index_buffer[2]), .ZN(n_1_0_2));
   NOR2_X1 i_1_0_15 (.A1(n_1_0_4), .A2(n_1_0_3), .ZN(n_12));
   NOR2_X1 i_1_0_16 (.A1(n_1_0_6), .A2(n_1_0_3), .ZN(n_13));
   NAND2_X1 i_1_0_17 (.A1(n_1_0_12), .A2(index_buffer[2]), .ZN(n_1_0_3));
   NOR2_X1 i_1_0_18 (.A1(n_1_0_5), .A2(n_1_0_4), .ZN(n_14));
   NAND3_X1 i_1_0_19 (.A1(index_buffer[3]), .A2(n_1_0_7), .A3(n_1_0_11), 
      .ZN(n_1_0_4));
   NOR2_X1 i_1_0_20 (.A1(n_1_0_6), .A2(n_1_0_5), .ZN(n_15));
   NAND2_X1 i_1_0_21 (.A1(index_buffer[2]), .A2(index_buffer[1]), .ZN(n_1_0_5));
   NAND3_X1 i_1_0_22 (.A1(index_buffer[3]), .A2(index_buffer[0]), .A3(n_1_0_7), 
      .ZN(n_1_0_6));
   AND4_X1 i_1_0_23 (.A1(bias_or_filter), .A2(n_1_0_8), .A3(n_1_0_14), .A4(
      n_1_0_10), .ZN(n_1_0_7));
   NOR4_X1 i_1_0_24 (.A1(n_1_0_9), .A2(index_buffer[5]), .A3(index_buffer[6]), 
      .A4(index_buffer[7]), .ZN(n_1_0_8));
   OR4_X1 i_1_0_25 (.A1(index_buffer[10]), .A2(index_buffer[9]), .A3(
      index_buffer[8]), .A4(index_buffer[4]), .ZN(n_1_0_9));
   NOR4_X1 i_1_0_26 (.A1(index_buffer[14]), .A2(index_buffer[13]), .A3(
      index_buffer[12]), .A4(index_buffer[11]), .ZN(n_1_0_10));
   INV_X1 i_1_0_27 (.A(index_buffer[0]), .ZN(n_1_0_11));
   INV_X1 i_1_0_28 (.A(index_buffer[1]), .ZN(n_1_0_12));
   INV_X1 i_1_0_29 (.A(index_buffer[3]), .ZN(n_1_0_13));
   INV_X1 i_1_0_30 (.A(index_buffer[15]), .ZN(n_1_0_14));
   NAND4_X1 i_2_44_0 (.A1(n_2_44_8), .A2(n_2_44_6), .A3(n_2_44_4), .A4(n_2_44_0), 
      .ZN(\output_filter[4][4] [0]));
   AOI221_X1 i_2_44_1 (.A(n_2_44_1), .B1(n_25), .B2(\buffer[0][4][4] [0]), 
      .C1(\buffer[12][4][4] [0]), .C2(n_27), .ZN(n_2_44_0));
   NAND4_X1 i_2_44_2 (.A1(n_2_44_7), .A2(n_2_44_5), .A3(n_2_44_3), .A4(n_2_44_2), 
      .ZN(n_2_44_1));
   AOI22_X1 i_2_44_3 (.A1(\buffer[15][4][4] [0]), .A2(n_22), .B1(n_29), .B2(
      \buffer[7][4][4] [0]), .ZN(n_2_44_2));
   AOI22_X1 i_2_44_4 (.A1(\buffer[10][4][4] [0]), .A2(n_21), .B1(n_16), .B2(
      \buffer[8][4][4] [0]), .ZN(n_2_44_3));
   AOI22_X1 i_2_44_5 (.A1(\buffer[6][4][4] [0]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][4] [0]), .ZN(n_2_44_4));
   AOI22_X1 i_2_44_6 (.A1(\buffer[9][4][4] [0]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][4] [0]), .ZN(n_2_44_5));
   AOI22_X1 i_2_44_7 (.A1(\buffer[14][4][4] [0]), .A2(n_19), .B1(n_23), .B2(
      \buffer[1][4][4] [0]), .ZN(n_2_44_6));
   AOI22_X1 i_2_44_8 (.A1(\buffer[11][4][4] [0]), .A2(n_17), .B1(n_18), .B2(
      \buffer[5][4][4] [0]), .ZN(n_2_44_7));
   AOI22_X1 i_2_44_9 (.A1(\buffer[13][4][4] [0]), .A2(n_26), .B1(n_24), .B2(
      \buffer[2][4][4] [0]), .ZN(n_2_44_8));
   NAND4_X1 i_2_44_10 (.A1(n_2_44_17), .A2(n_2_44_15), .A3(n_2_44_13), .A4(
      n_2_44_9), .ZN(\output_filter[4][4] [1]));
   AOI221_X1 i_2_44_11 (.A(n_2_44_10), .B1(n_25), .B2(\buffer[0][4][4] [1]), 
      .C1(\buffer[12][4][4] [1]), .C2(n_27), .ZN(n_2_44_9));
   NAND4_X1 i_2_44_12 (.A1(n_2_44_16), .A2(n_2_44_14), .A3(n_2_44_12), .A4(
      n_2_44_11), .ZN(n_2_44_10));
   AOI22_X1 i_2_44_13 (.A1(\buffer[15][4][4] [1]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][4] [1]), .ZN(n_2_44_11));
   AOI22_X1 i_2_44_14 (.A1(\buffer[10][4][4] [1]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][4] [1]), .ZN(n_2_44_12));
   AOI22_X1 i_2_44_15 (.A1(\buffer[6][4][4] [1]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][4] [1]), .ZN(n_2_44_13));
   AOI22_X1 i_2_44_16 (.A1(\buffer[9][4][4] [1]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][4] [1]), .ZN(n_2_44_14));
   AOI22_X1 i_2_44_17 (.A1(\buffer[14][4][4] [1]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][4] [1]), .ZN(n_2_44_15));
   AOI22_X1 i_2_44_18 (.A1(\buffer[11][4][4] [1]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][4] [1]), .ZN(n_2_44_16));
   AOI22_X1 i_2_44_19 (.A1(\buffer[13][4][4] [1]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][4] [1]), .ZN(n_2_44_17));
   NAND4_X1 i_2_44_20 (.A1(n_2_44_26), .A2(n_2_44_24), .A3(n_2_44_22), .A4(
      n_2_44_18), .ZN(\output_filter[4][4] [2]));
   AOI221_X1 i_2_44_21 (.A(n_2_44_19), .B1(n_25), .B2(\buffer[0][4][4] [2]), 
      .C1(\buffer[12][4][4] [2]), .C2(n_27), .ZN(n_2_44_18));
   NAND4_X1 i_2_44_22 (.A1(n_2_44_25), .A2(n_2_44_23), .A3(n_2_44_21), .A4(
      n_2_44_20), .ZN(n_2_44_19));
   AOI22_X1 i_2_44_23 (.A1(\buffer[15][4][4] [2]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][4] [2]), .ZN(n_2_44_20));
   AOI22_X1 i_2_44_24 (.A1(\buffer[10][4][4] [2]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][4] [2]), .ZN(n_2_44_21));
   AOI22_X1 i_2_44_25 (.A1(\buffer[6][4][4] [2]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][4] [2]), .ZN(n_2_44_22));
   AOI22_X1 i_2_44_26 (.A1(\buffer[9][4][4] [2]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][4] [2]), .ZN(n_2_44_23));
   AOI22_X1 i_2_44_27 (.A1(\buffer[14][4][4] [2]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][4] [2]), .ZN(n_2_44_24));
   AOI22_X1 i_2_44_28 (.A1(\buffer[11][4][4] [2]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][4] [2]), .ZN(n_2_44_25));
   AOI22_X1 i_2_44_29 (.A1(\buffer[13][4][4] [2]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][4] [2]), .ZN(n_2_44_26));
   NAND4_X1 i_2_44_30 (.A1(n_2_44_35), .A2(n_2_44_33), .A3(n_2_44_31), .A4(
      n_2_44_27), .ZN(\output_filter[4][4] [3]));
   AOI221_X1 i_2_44_31 (.A(n_2_44_28), .B1(n_25), .B2(\buffer[0][4][4] [3]), 
      .C1(\buffer[12][4][4] [3]), .C2(n_27), .ZN(n_2_44_27));
   NAND4_X1 i_2_44_32 (.A1(n_2_44_34), .A2(n_2_44_32), .A3(n_2_44_30), .A4(
      n_2_44_29), .ZN(n_2_44_28));
   AOI22_X1 i_2_44_33 (.A1(\buffer[15][4][4] [3]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][4] [3]), .ZN(n_2_44_29));
   AOI22_X1 i_2_44_34 (.A1(\buffer[10][4][4] [3]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][4] [3]), .ZN(n_2_44_30));
   AOI22_X1 i_2_44_35 (.A1(\buffer[6][4][4] [3]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][4] [3]), .ZN(n_2_44_31));
   AOI22_X1 i_2_44_36 (.A1(\buffer[9][4][4] [3]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][4] [3]), .ZN(n_2_44_32));
   AOI22_X1 i_2_44_37 (.A1(\buffer[14][4][4] [3]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][4] [3]), .ZN(n_2_44_33));
   AOI22_X1 i_2_44_38 (.A1(\buffer[11][4][4] [3]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][4] [3]), .ZN(n_2_44_34));
   AOI22_X1 i_2_44_39 (.A1(\buffer[13][4][4] [3]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][4] [3]), .ZN(n_2_44_35));
   NAND4_X1 i_2_44_40 (.A1(n_2_44_44), .A2(n_2_44_42), .A3(n_2_44_40), .A4(
      n_2_44_36), .ZN(\output_filter[4][4] [4]));
   AOI221_X1 i_2_44_41 (.A(n_2_44_37), .B1(n_25), .B2(\buffer[0][4][4] [4]), 
      .C1(\buffer[12][4][4] [4]), .C2(n_27), .ZN(n_2_44_36));
   NAND4_X1 i_2_44_42 (.A1(n_2_44_43), .A2(n_2_44_41), .A3(n_2_44_39), .A4(
      n_2_44_38), .ZN(n_2_44_37));
   AOI22_X1 i_2_44_43 (.A1(\buffer[15][4][4] [4]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][4] [4]), .ZN(n_2_44_38));
   AOI22_X1 i_2_44_44 (.A1(\buffer[10][4][4] [4]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][4] [4]), .ZN(n_2_44_39));
   AOI22_X1 i_2_44_45 (.A1(\buffer[6][4][4] [4]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][4] [4]), .ZN(n_2_44_40));
   AOI22_X1 i_2_44_46 (.A1(\buffer[9][4][4] [4]), .A2(n_20), .B1(n_24), .B2(
      \buffer[2][4][4] [4]), .ZN(n_2_44_41));
   AOI22_X1 i_2_44_47 (.A1(\buffer[14][4][4] [4]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][4] [4]), .ZN(n_2_44_42));
   AOI22_X1 i_2_44_48 (.A1(\buffer[11][4][4] [4]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][4] [4]), .ZN(n_2_44_43));
   AOI22_X1 i_2_44_49 (.A1(\buffer[13][4][4] [4]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][4][4] [4]), .ZN(n_2_44_44));
   NAND4_X1 i_2_44_50 (.A1(n_2_44_53), .A2(n_2_44_51), .A3(n_2_44_49), .A4(
      n_2_44_45), .ZN(\output_filter[4][4] [5]));
   AOI221_X1 i_2_44_51 (.A(n_2_44_46), .B1(n_25), .B2(\buffer[0][4][4] [5]), 
      .C1(\buffer[12][4][4] [5]), .C2(n_27), .ZN(n_2_44_45));
   NAND4_X1 i_2_44_52 (.A1(n_2_44_52), .A2(n_2_44_50), .A3(n_2_44_48), .A4(
      n_2_44_47), .ZN(n_2_44_46));
   AOI22_X1 i_2_44_53 (.A1(\buffer[15][4][4] [5]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][4] [5]), .ZN(n_2_44_47));
   AOI22_X1 i_2_44_54 (.A1(\buffer[10][4][4] [5]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][4] [5]), .ZN(n_2_44_48));
   AOI22_X1 i_2_44_55 (.A1(\buffer[6][4][4] [5]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][4] [5]), .ZN(n_2_44_49));
   AOI22_X1 i_2_44_56 (.A1(\buffer[9][4][4] [5]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][4] [5]), .ZN(n_2_44_50));
   AOI22_X1 i_2_44_57 (.A1(\buffer[14][4][4] [5]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][4] [5]), .ZN(n_2_44_51));
   AOI22_X1 i_2_44_58 (.A1(\buffer[11][4][4] [5]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][4] [5]), .ZN(n_2_44_52));
   AOI22_X1 i_2_44_59 (.A1(\buffer[13][4][4] [5]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][4] [5]), .ZN(n_2_44_53));
   NAND4_X1 i_2_44_60 (.A1(n_2_44_62), .A2(n_2_44_60), .A3(n_2_44_58), .A4(
      n_2_44_54), .ZN(\output_filter[4][4] [6]));
   AOI221_X1 i_2_44_61 (.A(n_2_44_55), .B1(n_25), .B2(\buffer[0][4][4] [6]), 
      .C1(\buffer[12][4][4] [6]), .C2(n_27), .ZN(n_2_44_54));
   NAND4_X1 i_2_44_62 (.A1(n_2_44_61), .A2(n_2_44_59), .A3(n_2_44_57), .A4(
      n_2_44_56), .ZN(n_2_44_55));
   AOI22_X1 i_2_44_63 (.A1(\buffer[15][4][4] [6]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][4] [6]), .ZN(n_2_44_56));
   AOI22_X1 i_2_44_64 (.A1(\buffer[10][4][4] [6]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][4] [6]), .ZN(n_2_44_57));
   AOI22_X1 i_2_44_65 (.A1(\buffer[6][4][4] [6]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][4] [6]), .ZN(n_2_44_58));
   AOI22_X1 i_2_44_66 (.A1(\buffer[9][4][4] [6]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][4] [6]), .ZN(n_2_44_59));
   AOI22_X1 i_2_44_67 (.A1(\buffer[14][4][4] [6]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][4] [6]), .ZN(n_2_44_60));
   AOI22_X1 i_2_44_68 (.A1(\buffer[11][4][4] [6]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][4] [6]), .ZN(n_2_44_61));
   AOI22_X1 i_2_44_69 (.A1(\buffer[13][4][4] [6]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][4] [6]), .ZN(n_2_44_62));
   NAND4_X1 i_2_44_70 (.A1(n_2_44_71), .A2(n_2_44_69), .A3(n_2_44_67), .A4(
      n_2_44_63), .ZN(\output_filter[4][4] [7]));
   AOI221_X1 i_2_44_71 (.A(n_2_44_64), .B1(n_25), .B2(\buffer[0][4][4] [7]), 
      .C1(\buffer[12][4][4] [7]), .C2(n_27), .ZN(n_2_44_63));
   NAND4_X1 i_2_44_72 (.A1(n_2_44_70), .A2(n_2_44_68), .A3(n_2_44_66), .A4(
      n_2_44_65), .ZN(n_2_44_64));
   AOI22_X1 i_2_44_73 (.A1(\buffer[15][4][4] [7]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][4] [7]), .ZN(n_2_44_65));
   AOI22_X1 i_2_44_74 (.A1(\buffer[10][4][4] [7]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][4] [7]), .ZN(n_2_44_66));
   AOI22_X1 i_2_44_75 (.A1(\buffer[6][4][4] [7]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][4] [7]), .ZN(n_2_44_67));
   AOI22_X1 i_2_44_76 (.A1(\buffer[9][4][4] [7]), .A2(n_20), .B1(n_24), .B2(
      \buffer[2][4][4] [7]), .ZN(n_2_44_68));
   AOI22_X1 i_2_44_77 (.A1(\buffer[14][4][4] [7]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][4] [7]), .ZN(n_2_44_69));
   AOI22_X1 i_2_44_78 (.A1(\buffer[11][4][4] [7]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][4] [7]), .ZN(n_2_44_70));
   AOI22_X1 i_2_44_79 (.A1(\buffer[13][4][4] [7]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][4][4] [7]), .ZN(n_2_44_71));
   NAND4_X1 i_2_44_80 (.A1(n_2_44_80), .A2(n_2_44_78), .A3(n_2_44_76), .A4(
      n_2_44_72), .ZN(\output_filter[4][4] [8]));
   AOI221_X1 i_2_44_81 (.A(n_2_44_73), .B1(n_25), .B2(\buffer[0][4][4] [8]), 
      .C1(\buffer[12][4][4] [8]), .C2(n_27), .ZN(n_2_44_72));
   NAND4_X1 i_2_44_82 (.A1(n_2_44_79), .A2(n_2_44_77), .A3(n_2_44_75), .A4(
      n_2_44_74), .ZN(n_2_44_73));
   AOI22_X1 i_2_44_83 (.A1(\buffer[15][4][4] [8]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][4] [8]), .ZN(n_2_44_74));
   AOI22_X1 i_2_44_84 (.A1(\buffer[10][4][4] [8]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][4] [8]), .ZN(n_2_44_75));
   AOI22_X1 i_2_44_85 (.A1(\buffer[6][4][4] [8]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][4] [8]), .ZN(n_2_44_76));
   AOI22_X1 i_2_44_86 (.A1(\buffer[9][4][4] [8]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][4] [8]), .ZN(n_2_44_77));
   AOI22_X1 i_2_44_87 (.A1(\buffer[14][4][4] [8]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][4] [8]), .ZN(n_2_44_78));
   AOI22_X1 i_2_44_88 (.A1(\buffer[11][4][4] [8]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][4] [8]), .ZN(n_2_44_79));
   AOI22_X1 i_2_44_89 (.A1(\buffer[13][4][4] [8]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][4] [8]), .ZN(n_2_44_80));
   NAND4_X1 i_2_44_90 (.A1(n_2_44_89), .A2(n_2_44_87), .A3(n_2_44_85), .A4(
      n_2_44_81), .ZN(\output_filter[4][4] [9]));
   AOI221_X1 i_2_44_91 (.A(n_2_44_82), .B1(n_25), .B2(\buffer[0][4][4] [9]), 
      .C1(\buffer[12][4][4] [9]), .C2(n_27), .ZN(n_2_44_81));
   NAND4_X1 i_2_44_92 (.A1(n_2_44_88), .A2(n_2_44_86), .A3(n_2_44_84), .A4(
      n_2_44_83), .ZN(n_2_44_82));
   AOI22_X1 i_2_44_93 (.A1(\buffer[15][4][4] [9]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][4] [9]), .ZN(n_2_44_83));
   AOI22_X1 i_2_44_94 (.A1(\buffer[10][4][4] [9]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][4] [9]), .ZN(n_2_44_84));
   AOI22_X1 i_2_44_95 (.A1(\buffer[6][4][4] [9]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][4] [9]), .ZN(n_2_44_85));
   AOI22_X1 i_2_44_96 (.A1(\buffer[9][4][4] [9]), .A2(n_20), .B1(n_24), .B2(
      \buffer[2][4][4] [9]), .ZN(n_2_44_86));
   AOI22_X1 i_2_44_97 (.A1(\buffer[14][4][4] [9]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][4] [9]), .ZN(n_2_44_87));
   AOI22_X1 i_2_44_98 (.A1(\buffer[11][4][4] [9]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][4] [9]), .ZN(n_2_44_88));
   AOI22_X1 i_2_44_99 (.A1(\buffer[13][4][4] [9]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][4][4] [9]), .ZN(n_2_44_89));
   NAND4_X1 i_2_44_100 (.A1(n_2_44_98), .A2(n_2_44_96), .A3(n_2_44_94), .A4(
      n_2_44_90), .ZN(\output_filter[4][4] [10]));
   AOI221_X1 i_2_44_101 (.A(n_2_44_91), .B1(n_25), .B2(\buffer[0][4][4] [10]), 
      .C1(\buffer[12][4][4] [10]), .C2(n_27), .ZN(n_2_44_90));
   NAND4_X1 i_2_44_102 (.A1(n_2_44_97), .A2(n_2_44_95), .A3(n_2_44_93), .A4(
      n_2_44_92), .ZN(n_2_44_91));
   AOI22_X1 i_2_44_103 (.A1(\buffer[15][4][4] [10]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][4] [10]), .ZN(n_2_44_92));
   AOI22_X1 i_2_44_104 (.A1(\buffer[10][4][4] [10]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][4] [10]), .ZN(n_2_44_93));
   AOI22_X1 i_2_44_105 (.A1(\buffer[6][4][4] [10]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][4][4] [10]), .ZN(n_2_44_94));
   AOI22_X1 i_2_44_106 (.A1(\buffer[9][4][4] [10]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][4][4] [10]), .ZN(n_2_44_95));
   AOI22_X1 i_2_44_107 (.A1(\buffer[14][4][4] [10]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][4] [10]), .ZN(n_2_44_96));
   AOI22_X1 i_2_44_108 (.A1(\buffer[11][4][4] [10]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][4] [10]), .ZN(n_2_44_97));
   AOI22_X1 i_2_44_109 (.A1(\buffer[13][4][4] [10]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][4] [10]), .ZN(n_2_44_98));
   NAND4_X1 i_2_44_110 (.A1(n_2_44_107), .A2(n_2_44_105), .A3(n_2_44_103), 
      .A4(n_2_44_99), .ZN(\output_filter[4][4] [11]));
   AOI221_X1 i_2_44_111 (.A(n_2_44_100), .B1(n_25), .B2(\buffer[0][4][4] [11]), 
      .C1(\buffer[12][4][4] [11]), .C2(n_27), .ZN(n_2_44_99));
   NAND4_X1 i_2_44_112 (.A1(n_2_44_106), .A2(n_2_44_104), .A3(n_2_44_102), 
      .A4(n_2_44_101), .ZN(n_2_44_100));
   AOI22_X1 i_2_44_113 (.A1(\buffer[15][4][4] [11]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][4] [11]), .ZN(n_2_44_101));
   AOI22_X1 i_2_44_114 (.A1(\buffer[10][4][4] [11]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][4] [11]), .ZN(n_2_44_102));
   AOI22_X1 i_2_44_115 (.A1(\buffer[6][4][4] [11]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][4][4] [11]), .ZN(n_2_44_103));
   AOI22_X1 i_2_44_116 (.A1(\buffer[9][4][4] [11]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][4][4] [11]), .ZN(n_2_44_104));
   AOI22_X1 i_2_44_117 (.A1(\buffer[14][4][4] [11]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][4] [11]), .ZN(n_2_44_105));
   AOI22_X1 i_2_44_118 (.A1(\buffer[11][4][4] [11]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][4] [11]), .ZN(n_2_44_106));
   AOI22_X1 i_2_44_119 (.A1(\buffer[13][4][4] [11]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][4][4] [11]), .ZN(n_2_44_107));
   NAND4_X1 i_2_44_120 (.A1(n_2_44_116), .A2(n_2_44_114), .A3(n_2_44_112), 
      .A4(n_2_44_108), .ZN(\output_filter[4][4] [12]));
   AOI221_X1 i_2_44_121 (.A(n_2_44_109), .B1(n_25), .B2(\buffer[0][4][4] [12]), 
      .C1(\buffer[12][4][4] [12]), .C2(n_27), .ZN(n_2_44_108));
   NAND4_X1 i_2_44_122 (.A1(n_2_44_115), .A2(n_2_44_113), .A3(n_2_44_111), 
      .A4(n_2_44_110), .ZN(n_2_44_109));
   AOI22_X1 i_2_44_123 (.A1(\buffer[15][4][4] [12]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][4] [12]), .ZN(n_2_44_110));
   AOI22_X1 i_2_44_124 (.A1(\buffer[10][4][4] [12]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][4] [12]), .ZN(n_2_44_111));
   AOI22_X1 i_2_44_125 (.A1(\buffer[6][4][4] [12]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][4][4] [12]), .ZN(n_2_44_112));
   AOI22_X1 i_2_44_126 (.A1(\buffer[9][4][4] [12]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][4][4] [12]), .ZN(n_2_44_113));
   AOI22_X1 i_2_44_127 (.A1(\buffer[14][4][4] [12]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][4] [12]), .ZN(n_2_44_114));
   AOI22_X1 i_2_44_128 (.A1(\buffer[11][4][4] [12]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][4] [12]), .ZN(n_2_44_115));
   AOI22_X1 i_2_44_129 (.A1(\buffer[13][4][4] [12]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][4] [12]), .ZN(n_2_44_116));
   NAND4_X1 i_2_44_130 (.A1(n_2_44_125), .A2(n_2_44_123), .A3(n_2_44_121), 
      .A4(n_2_44_117), .ZN(\output_filter[4][4] [13]));
   AOI221_X1 i_2_44_131 (.A(n_2_44_118), .B1(n_25), .B2(\buffer[0][4][4] [13]), 
      .C1(\buffer[12][4][4] [13]), .C2(n_27), .ZN(n_2_44_117));
   NAND4_X1 i_2_44_132 (.A1(n_2_44_124), .A2(n_2_44_122), .A3(n_2_44_120), 
      .A4(n_2_44_119), .ZN(n_2_44_118));
   AOI22_X1 i_2_44_133 (.A1(\buffer[15][4][4] [13]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][4] [13]), .ZN(n_2_44_119));
   AOI22_X1 i_2_44_134 (.A1(\buffer[10][4][4] [13]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][4] [13]), .ZN(n_2_44_120));
   AOI22_X1 i_2_44_135 (.A1(\buffer[6][4][4] [13]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][4][4] [13]), .ZN(n_2_44_121));
   AOI22_X1 i_2_44_136 (.A1(\buffer[9][4][4] [13]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][4][4] [13]), .ZN(n_2_44_122));
   AOI22_X1 i_2_44_137 (.A1(\buffer[14][4][4] [13]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][4] [13]), .ZN(n_2_44_123));
   AOI22_X1 i_2_44_138 (.A1(\buffer[11][4][4] [13]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][4] [13]), .ZN(n_2_44_124));
   AOI22_X1 i_2_44_139 (.A1(\buffer[13][4][4] [13]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][4][4] [13]), .ZN(n_2_44_125));
   NAND4_X1 i_2_44_140 (.A1(n_2_44_134), .A2(n_2_44_132), .A3(n_2_44_130), 
      .A4(n_2_44_126), .ZN(\output_filter[4][4] [14]));
   AOI221_X1 i_2_44_141 (.A(n_2_44_127), .B1(n_25), .B2(\buffer[0][4][4] [14]), 
      .C1(\buffer[12][4][4] [14]), .C2(n_27), .ZN(n_2_44_126));
   NAND4_X1 i_2_44_142 (.A1(n_2_44_133), .A2(n_2_44_131), .A3(n_2_44_129), 
      .A4(n_2_44_128), .ZN(n_2_44_127));
   AOI22_X1 i_2_44_143 (.A1(\buffer[15][4][4] [14]), .A2(n_22), .B1(n_16), 
      .B2(\buffer[8][4][4] [14]), .ZN(n_2_44_128));
   AOI22_X1 i_2_44_144 (.A1(\buffer[10][4][4] [14]), .A2(n_21), .B1(n_29), 
      .B2(\buffer[7][4][4] [14]), .ZN(n_2_44_129));
   AOI22_X1 i_2_44_145 (.A1(\buffer[6][4][4] [14]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][4][4] [14]), .ZN(n_2_44_130));
   AOI22_X1 i_2_44_146 (.A1(\buffer[9][4][4] [14]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][4][4] [14]), .ZN(n_2_44_131));
   AOI22_X1 i_2_44_147 (.A1(\buffer[14][4][4] [14]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][4] [14]), .ZN(n_2_44_132));
   AOI22_X1 i_2_44_148 (.A1(\buffer[11][4][4] [14]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][4] [14]), .ZN(n_2_44_133));
   AOI22_X1 i_2_44_149 (.A1(\buffer[13][4][4] [14]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][4] [14]), .ZN(n_2_44_134));
   NAND2_X1 i_2_44_150 (.A1(n_2_44_137), .A2(n_2_44_135), .ZN(
      \output_filter[4][4] [15]));
   AOI221_X1 i_2_44_151 (.A(n_2_44_136), .B1(n_31), .B2(\buffer[3][4][4] [15]), 
      .C1(\buffer[14][4][4] [15]), .C2(n_19), .ZN(n_2_44_135));
   NAND3_X1 i_2_44_152 (.A1(n_2_44_143), .A2(n_2_44_141), .A3(n_2_44_139), 
      .ZN(n_2_44_136));
   AOI221_X1 i_2_44_153 (.A(n_2_44_138), .B1(n_16), .B2(\buffer[8][4][4] [15]), 
      .C1(\buffer[13][4][4] [15]), .C2(n_26), .ZN(n_2_44_137));
   NAND3_X1 i_2_44_154 (.A1(n_2_44_144), .A2(n_2_44_142), .A3(n_2_44_140), 
      .ZN(n_2_44_138));
   AOI22_X1 i_2_44_155 (.A1(\buffer[11][4][4] [15]), .A2(n_17), .B1(n_24), 
      .B2(\buffer[2][4][4] [15]), .ZN(n_2_44_139));
   AOI22_X1 i_2_44_156 (.A1(\buffer[10][4][4] [15]), .A2(n_21), .B1(n_23), 
      .B2(\buffer[1][4][4] [15]), .ZN(n_2_44_140));
   AOI22_X1 i_2_44_157 (.A1(\buffer[6][4][4] [15]), .A2(n_28), .B1(n_18), 
      .B2(\buffer[5][4][4] [15]), .ZN(n_2_44_141));
   AOI22_X1 i_2_44_158 (.A1(\buffer[9][4][4] [15]), .A2(n_20), .B1(n_30), 
      .B2(\buffer[4][4][4] [15]), .ZN(n_2_44_142));
   AOI22_X1 i_2_44_159 (.A1(\buffer[7][4][4] [15]), .A2(n_29), .B1(n_25), 
      .B2(\buffer[0][4][4] [15]), .ZN(n_2_44_143));
   AOI22_X1 i_2_44_160 (.A1(\buffer[15][4][4] [15]), .A2(n_22), .B1(n_27), 
      .B2(\buffer[12][4][4] [15]), .ZN(n_2_44_144));
   NAND4_X1 i_3_43_0 (.A1(n_3_43_8), .A2(n_3_43_6), .A3(n_3_43_4), .A4(n_3_43_0), 
      .ZN(\output_filter[4][3] [0]));
   AOI221_X1 i_3_43_1 (.A(n_3_43_1), .B1(n_25), .B2(\buffer[0][4][3] [0]), 
      .C1(\buffer[12][4][3] [0]), .C2(n_27), .ZN(n_3_43_0));
   NAND4_X1 i_3_43_2 (.A1(n_3_43_7), .A2(n_3_43_5), .A3(n_3_43_3), .A4(n_3_43_2), 
      .ZN(n_3_43_1));
   AOI22_X1 i_3_43_3 (.A1(\buffer[15][4][3] [0]), .A2(n_22), .B1(n_29), .B2(
      \buffer[7][4][3] [0]), .ZN(n_3_43_2));
   AOI22_X1 i_3_43_4 (.A1(\buffer[10][4][3] [0]), .A2(n_21), .B1(n_16), .B2(
      \buffer[8][4][3] [0]), .ZN(n_3_43_3));
   AOI22_X1 i_3_43_5 (.A1(\buffer[6][4][3] [0]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][3] [0]), .ZN(n_3_43_4));
   AOI22_X1 i_3_43_6 (.A1(\buffer[9][4][3] [0]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][3] [0]), .ZN(n_3_43_5));
   AOI22_X1 i_3_43_7 (.A1(\buffer[14][4][3] [0]), .A2(n_19), .B1(n_23), .B2(
      \buffer[1][4][3] [0]), .ZN(n_3_43_6));
   AOI22_X1 i_3_43_8 (.A1(\buffer[11][4][3] [0]), .A2(n_17), .B1(n_18), .B2(
      \buffer[5][4][3] [0]), .ZN(n_3_43_7));
   AOI22_X1 i_3_43_9 (.A1(\buffer[13][4][3] [0]), .A2(n_26), .B1(n_24), .B2(
      \buffer[2][4][3] [0]), .ZN(n_3_43_8));
   NAND4_X1 i_3_43_10 (.A1(n_3_43_17), .A2(n_3_43_15), .A3(n_3_43_13), .A4(
      n_3_43_9), .ZN(\output_filter[4][3] [1]));
   AOI221_X1 i_3_43_11 (.A(n_3_43_10), .B1(n_25), .B2(\buffer[0][4][3] [1]), 
      .C1(\buffer[12][4][3] [1]), .C2(n_27), .ZN(n_3_43_9));
   NAND4_X1 i_3_43_12 (.A1(n_3_43_16), .A2(n_3_43_14), .A3(n_3_43_12), .A4(
      n_3_43_11), .ZN(n_3_43_10));
   AOI22_X1 i_3_43_13 (.A1(\buffer[15][4][3] [1]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][3] [1]), .ZN(n_3_43_11));
   AOI22_X1 i_3_43_14 (.A1(\buffer[10][4][3] [1]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][3] [1]), .ZN(n_3_43_12));
   AOI22_X1 i_3_43_15 (.A1(\buffer[6][4][3] [1]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][3] [1]), .ZN(n_3_43_13));
   AOI22_X1 i_3_43_16 (.A1(\buffer[9][4][3] [1]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][3] [1]), .ZN(n_3_43_14));
   AOI22_X1 i_3_43_17 (.A1(\buffer[14][4][3] [1]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][3] [1]), .ZN(n_3_43_15));
   AOI22_X1 i_3_43_18 (.A1(\buffer[11][4][3] [1]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][3] [1]), .ZN(n_3_43_16));
   AOI22_X1 i_3_43_19 (.A1(\buffer[13][4][3] [1]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][3] [1]), .ZN(n_3_43_17));
   NAND4_X1 i_3_43_20 (.A1(n_3_43_26), .A2(n_3_43_24), .A3(n_3_43_22), .A4(
      n_3_43_18), .ZN(\output_filter[4][3] [2]));
   AOI221_X1 i_3_43_21 (.A(n_3_43_19), .B1(n_25), .B2(\buffer[0][4][3] [2]), 
      .C1(\buffer[12][4][3] [2]), .C2(n_27), .ZN(n_3_43_18));
   NAND4_X1 i_3_43_22 (.A1(n_3_43_25), .A2(n_3_43_23), .A3(n_3_43_21), .A4(
      n_3_43_20), .ZN(n_3_43_19));
   AOI22_X1 i_3_43_23 (.A1(\buffer[15][4][3] [2]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][3] [2]), .ZN(n_3_43_20));
   AOI22_X1 i_3_43_24 (.A1(\buffer[10][4][3] [2]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][3] [2]), .ZN(n_3_43_21));
   AOI22_X1 i_3_43_25 (.A1(\buffer[6][4][3] [2]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][3] [2]), .ZN(n_3_43_22));
   AOI22_X1 i_3_43_26 (.A1(\buffer[9][4][3] [2]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][3] [2]), .ZN(n_3_43_23));
   AOI22_X1 i_3_43_27 (.A1(\buffer[14][4][3] [2]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][3] [2]), .ZN(n_3_43_24));
   AOI22_X1 i_3_43_28 (.A1(\buffer[11][4][3] [2]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][3] [2]), .ZN(n_3_43_25));
   AOI22_X1 i_3_43_29 (.A1(\buffer[13][4][3] [2]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][3] [2]), .ZN(n_3_43_26));
   NAND4_X1 i_3_43_30 (.A1(n_3_43_35), .A2(n_3_43_33), .A3(n_3_43_31), .A4(
      n_3_43_27), .ZN(\output_filter[4][3] [3]));
   AOI221_X1 i_3_43_31 (.A(n_3_43_28), .B1(n_25), .B2(\buffer[0][4][3] [3]), 
      .C1(\buffer[12][4][3] [3]), .C2(n_27), .ZN(n_3_43_27));
   NAND4_X1 i_3_43_32 (.A1(n_3_43_34), .A2(n_3_43_32), .A3(n_3_43_30), .A4(
      n_3_43_29), .ZN(n_3_43_28));
   AOI22_X1 i_3_43_33 (.A1(\buffer[15][4][3] [3]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][3] [3]), .ZN(n_3_43_29));
   AOI22_X1 i_3_43_34 (.A1(\buffer[10][4][3] [3]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][3] [3]), .ZN(n_3_43_30));
   AOI22_X1 i_3_43_35 (.A1(\buffer[6][4][3] [3]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][3] [3]), .ZN(n_3_43_31));
   AOI22_X1 i_3_43_36 (.A1(\buffer[9][4][3] [3]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][3] [3]), .ZN(n_3_43_32));
   AOI22_X1 i_3_43_37 (.A1(\buffer[14][4][3] [3]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][3] [3]), .ZN(n_3_43_33));
   AOI22_X1 i_3_43_38 (.A1(\buffer[11][4][3] [3]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][3] [3]), .ZN(n_3_43_34));
   AOI22_X1 i_3_43_39 (.A1(\buffer[13][4][3] [3]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][3] [3]), .ZN(n_3_43_35));
   NAND4_X1 i_3_43_40 (.A1(n_3_43_44), .A2(n_3_43_42), .A3(n_3_43_40), .A4(
      n_3_43_36), .ZN(\output_filter[4][3] [4]));
   AOI221_X1 i_3_43_41 (.A(n_3_43_37), .B1(n_25), .B2(\buffer[0][4][3] [4]), 
      .C1(\buffer[12][4][3] [4]), .C2(n_27), .ZN(n_3_43_36));
   NAND4_X1 i_3_43_42 (.A1(n_3_43_43), .A2(n_3_43_41), .A3(n_3_43_39), .A4(
      n_3_43_38), .ZN(n_3_43_37));
   AOI22_X1 i_3_43_43 (.A1(\buffer[15][4][3] [4]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][3] [4]), .ZN(n_3_43_38));
   AOI22_X1 i_3_43_44 (.A1(\buffer[10][4][3] [4]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][3] [4]), .ZN(n_3_43_39));
   AOI22_X1 i_3_43_45 (.A1(\buffer[6][4][3] [4]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][3] [4]), .ZN(n_3_43_40));
   AOI22_X1 i_3_43_46 (.A1(\buffer[9][4][3] [4]), .A2(n_20), .B1(n_24), .B2(
      \buffer[2][4][3] [4]), .ZN(n_3_43_41));
   AOI22_X1 i_3_43_47 (.A1(\buffer[14][4][3] [4]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][3] [4]), .ZN(n_3_43_42));
   AOI22_X1 i_3_43_48 (.A1(\buffer[11][4][3] [4]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][3] [4]), .ZN(n_3_43_43));
   AOI22_X1 i_3_43_49 (.A1(\buffer[13][4][3] [4]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][4][3] [4]), .ZN(n_3_43_44));
   NAND4_X1 i_3_43_50 (.A1(n_3_43_53), .A2(n_3_43_51), .A3(n_3_43_49), .A4(
      n_3_43_45), .ZN(\output_filter[4][3] [5]));
   AOI221_X1 i_3_43_51 (.A(n_3_43_46), .B1(n_25), .B2(\buffer[0][4][3] [5]), 
      .C1(\buffer[12][4][3] [5]), .C2(n_27), .ZN(n_3_43_45));
   NAND4_X1 i_3_43_52 (.A1(n_3_43_52), .A2(n_3_43_50), .A3(n_3_43_48), .A4(
      n_3_43_47), .ZN(n_3_43_46));
   AOI22_X1 i_3_43_53 (.A1(\buffer[15][4][3] [5]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][3] [5]), .ZN(n_3_43_47));
   AOI22_X1 i_3_43_54 (.A1(\buffer[10][4][3] [5]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][3] [5]), .ZN(n_3_43_48));
   AOI22_X1 i_3_43_55 (.A1(\buffer[6][4][3] [5]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][3] [5]), .ZN(n_3_43_49));
   AOI22_X1 i_3_43_56 (.A1(\buffer[9][4][3] [5]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][3] [5]), .ZN(n_3_43_50));
   AOI22_X1 i_3_43_57 (.A1(\buffer[14][4][3] [5]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][3] [5]), .ZN(n_3_43_51));
   AOI22_X1 i_3_43_58 (.A1(\buffer[11][4][3] [5]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][3] [5]), .ZN(n_3_43_52));
   AOI22_X1 i_3_43_59 (.A1(\buffer[13][4][3] [5]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][3] [5]), .ZN(n_3_43_53));
   NAND4_X1 i_3_43_60 (.A1(n_3_43_62), .A2(n_3_43_60), .A3(n_3_43_58), .A4(
      n_3_43_54), .ZN(\output_filter[4][3] [6]));
   AOI221_X1 i_3_43_61 (.A(n_3_43_55), .B1(n_25), .B2(\buffer[0][4][3] [6]), 
      .C1(\buffer[12][4][3] [6]), .C2(n_27), .ZN(n_3_43_54));
   NAND4_X1 i_3_43_62 (.A1(n_3_43_61), .A2(n_3_43_59), .A3(n_3_43_57), .A4(
      n_3_43_56), .ZN(n_3_43_55));
   AOI22_X1 i_3_43_63 (.A1(\buffer[15][4][3] [6]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][3] [6]), .ZN(n_3_43_56));
   AOI22_X1 i_3_43_64 (.A1(\buffer[10][4][3] [6]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][3] [6]), .ZN(n_3_43_57));
   AOI22_X1 i_3_43_65 (.A1(\buffer[6][4][3] [6]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][3] [6]), .ZN(n_3_43_58));
   AOI22_X1 i_3_43_66 (.A1(\buffer[9][4][3] [6]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][3] [6]), .ZN(n_3_43_59));
   AOI22_X1 i_3_43_67 (.A1(\buffer[14][4][3] [6]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][3] [6]), .ZN(n_3_43_60));
   AOI22_X1 i_3_43_68 (.A1(\buffer[11][4][3] [6]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][3] [6]), .ZN(n_3_43_61));
   AOI22_X1 i_3_43_69 (.A1(\buffer[13][4][3] [6]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][3] [6]), .ZN(n_3_43_62));
   NAND4_X1 i_3_43_70 (.A1(n_3_43_71), .A2(n_3_43_69), .A3(n_3_43_67), .A4(
      n_3_43_63), .ZN(\output_filter[4][3] [7]));
   AOI221_X1 i_3_43_71 (.A(n_3_43_64), .B1(n_25), .B2(\buffer[0][4][3] [7]), 
      .C1(\buffer[12][4][3] [7]), .C2(n_27), .ZN(n_3_43_63));
   NAND4_X1 i_3_43_72 (.A1(n_3_43_70), .A2(n_3_43_68), .A3(n_3_43_66), .A4(
      n_3_43_65), .ZN(n_3_43_64));
   AOI22_X1 i_3_43_73 (.A1(\buffer[15][4][3] [7]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][3] [7]), .ZN(n_3_43_65));
   AOI22_X1 i_3_43_74 (.A1(\buffer[10][4][3] [7]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][3] [7]), .ZN(n_3_43_66));
   AOI22_X1 i_3_43_75 (.A1(\buffer[6][4][3] [7]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][3] [7]), .ZN(n_3_43_67));
   AOI22_X1 i_3_43_76 (.A1(\buffer[9][4][3] [7]), .A2(n_20), .B1(n_24), .B2(
      \buffer[2][4][3] [7]), .ZN(n_3_43_68));
   AOI22_X1 i_3_43_77 (.A1(\buffer[14][4][3] [7]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][3] [7]), .ZN(n_3_43_69));
   AOI22_X1 i_3_43_78 (.A1(\buffer[11][4][3] [7]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][3] [7]), .ZN(n_3_43_70));
   AOI22_X1 i_3_43_79 (.A1(\buffer[13][4][3] [7]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][4][3] [7]), .ZN(n_3_43_71));
   NAND4_X1 i_3_43_80 (.A1(n_3_43_80), .A2(n_3_43_78), .A3(n_3_43_76), .A4(
      n_3_43_72), .ZN(\output_filter[4][3] [8]));
   AOI221_X1 i_3_43_81 (.A(n_3_43_73), .B1(n_25), .B2(\buffer[0][4][3] [8]), 
      .C1(\buffer[12][4][3] [8]), .C2(n_27), .ZN(n_3_43_72));
   NAND4_X1 i_3_43_82 (.A1(n_3_43_79), .A2(n_3_43_77), .A3(n_3_43_75), .A4(
      n_3_43_74), .ZN(n_3_43_73));
   AOI22_X1 i_3_43_83 (.A1(\buffer[15][4][3] [8]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][3] [8]), .ZN(n_3_43_74));
   AOI22_X1 i_3_43_84 (.A1(\buffer[10][4][3] [8]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][3] [8]), .ZN(n_3_43_75));
   AOI22_X1 i_3_43_85 (.A1(\buffer[6][4][3] [8]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][3] [8]), .ZN(n_3_43_76));
   AOI22_X1 i_3_43_86 (.A1(\buffer[9][4][3] [8]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][3] [8]), .ZN(n_3_43_77));
   AOI22_X1 i_3_43_87 (.A1(\buffer[14][4][3] [8]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][3] [8]), .ZN(n_3_43_78));
   AOI22_X1 i_3_43_88 (.A1(\buffer[11][4][3] [8]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][3] [8]), .ZN(n_3_43_79));
   AOI22_X1 i_3_43_89 (.A1(\buffer[13][4][3] [8]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][3] [8]), .ZN(n_3_43_80));
   NAND4_X1 i_3_43_90 (.A1(n_3_43_89), .A2(n_3_43_87), .A3(n_3_43_85), .A4(
      n_3_43_81), .ZN(\output_filter[4][3] [9]));
   AOI221_X1 i_3_43_91 (.A(n_3_43_82), .B1(n_25), .B2(\buffer[0][4][3] [9]), 
      .C1(\buffer[12][4][3] [9]), .C2(n_27), .ZN(n_3_43_81));
   NAND4_X1 i_3_43_92 (.A1(n_3_43_88), .A2(n_3_43_86), .A3(n_3_43_84), .A4(
      n_3_43_83), .ZN(n_3_43_82));
   AOI22_X1 i_3_43_93 (.A1(\buffer[15][4][3] [9]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][3] [9]), .ZN(n_3_43_83));
   AOI22_X1 i_3_43_94 (.A1(\buffer[10][4][3] [9]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][3] [9]), .ZN(n_3_43_84));
   AOI22_X1 i_3_43_95 (.A1(\buffer[6][4][3] [9]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][3] [9]), .ZN(n_3_43_85));
   AOI22_X1 i_3_43_96 (.A1(\buffer[9][4][3] [9]), .A2(n_20), .B1(n_24), .B2(
      \buffer[2][4][3] [9]), .ZN(n_3_43_86));
   AOI22_X1 i_3_43_97 (.A1(\buffer[14][4][3] [9]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][3] [9]), .ZN(n_3_43_87));
   AOI22_X1 i_3_43_98 (.A1(\buffer[11][4][3] [9]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][3] [9]), .ZN(n_3_43_88));
   AOI22_X1 i_3_43_99 (.A1(\buffer[13][4][3] [9]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][4][3] [9]), .ZN(n_3_43_89));
   NAND4_X1 i_3_43_100 (.A1(n_3_43_98), .A2(n_3_43_96), .A3(n_3_43_94), .A4(
      n_3_43_90), .ZN(\output_filter[4][3] [10]));
   AOI221_X1 i_3_43_101 (.A(n_3_43_91), .B1(n_25), .B2(\buffer[0][4][3] [10]), 
      .C1(\buffer[12][4][3] [10]), .C2(n_27), .ZN(n_3_43_90));
   NAND4_X1 i_3_43_102 (.A1(n_3_43_97), .A2(n_3_43_95), .A3(n_3_43_93), .A4(
      n_3_43_92), .ZN(n_3_43_91));
   AOI22_X1 i_3_43_103 (.A1(\buffer[15][4][3] [10]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][3] [10]), .ZN(n_3_43_92));
   AOI22_X1 i_3_43_104 (.A1(\buffer[10][4][3] [10]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][3] [10]), .ZN(n_3_43_93));
   AOI22_X1 i_3_43_105 (.A1(\buffer[6][4][3] [10]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][4][3] [10]), .ZN(n_3_43_94));
   AOI22_X1 i_3_43_106 (.A1(\buffer[9][4][3] [10]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][4][3] [10]), .ZN(n_3_43_95));
   AOI22_X1 i_3_43_107 (.A1(\buffer[14][4][3] [10]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][3] [10]), .ZN(n_3_43_96));
   AOI22_X1 i_3_43_108 (.A1(\buffer[11][4][3] [10]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][3] [10]), .ZN(n_3_43_97));
   AOI22_X1 i_3_43_109 (.A1(\buffer[13][4][3] [10]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][3] [10]), .ZN(n_3_43_98));
   NAND4_X1 i_3_43_110 (.A1(n_3_43_107), .A2(n_3_43_105), .A3(n_3_43_103), 
      .A4(n_3_43_99), .ZN(\output_filter[4][3] [11]));
   AOI221_X1 i_3_43_111 (.A(n_3_43_100), .B1(n_25), .B2(\buffer[0][4][3] [11]), 
      .C1(\buffer[12][4][3] [11]), .C2(n_27), .ZN(n_3_43_99));
   NAND4_X1 i_3_43_112 (.A1(n_3_43_106), .A2(n_3_43_104), .A3(n_3_43_102), 
      .A4(n_3_43_101), .ZN(n_3_43_100));
   AOI22_X1 i_3_43_113 (.A1(\buffer[15][4][3] [11]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][3] [11]), .ZN(n_3_43_101));
   AOI22_X1 i_3_43_114 (.A1(\buffer[10][4][3] [11]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][3] [11]), .ZN(n_3_43_102));
   AOI22_X1 i_3_43_115 (.A1(\buffer[6][4][3] [11]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][4][3] [11]), .ZN(n_3_43_103));
   AOI22_X1 i_3_43_116 (.A1(\buffer[9][4][3] [11]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][4][3] [11]), .ZN(n_3_43_104));
   AOI22_X1 i_3_43_117 (.A1(\buffer[14][4][3] [11]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][3] [11]), .ZN(n_3_43_105));
   AOI22_X1 i_3_43_118 (.A1(\buffer[11][4][3] [11]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][3] [11]), .ZN(n_3_43_106));
   AOI22_X1 i_3_43_119 (.A1(\buffer[13][4][3] [11]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][4][3] [11]), .ZN(n_3_43_107));
   NAND4_X1 i_3_43_120 (.A1(n_3_43_116), .A2(n_3_43_114), .A3(n_3_43_112), 
      .A4(n_3_43_108), .ZN(\output_filter[4][3] [12]));
   AOI221_X1 i_3_43_121 (.A(n_3_43_109), .B1(n_25), .B2(\buffer[0][4][3] [12]), 
      .C1(\buffer[12][4][3] [12]), .C2(n_27), .ZN(n_3_43_108));
   NAND4_X1 i_3_43_122 (.A1(n_3_43_115), .A2(n_3_43_113), .A3(n_3_43_111), 
      .A4(n_3_43_110), .ZN(n_3_43_109));
   AOI22_X1 i_3_43_123 (.A1(\buffer[15][4][3] [12]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][3] [12]), .ZN(n_3_43_110));
   AOI22_X1 i_3_43_124 (.A1(\buffer[10][4][3] [12]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][3] [12]), .ZN(n_3_43_111));
   AOI22_X1 i_3_43_125 (.A1(\buffer[6][4][3] [12]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][4][3] [12]), .ZN(n_3_43_112));
   AOI22_X1 i_3_43_126 (.A1(\buffer[9][4][3] [12]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][4][3] [12]), .ZN(n_3_43_113));
   AOI22_X1 i_3_43_127 (.A1(\buffer[14][4][3] [12]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][3] [12]), .ZN(n_3_43_114));
   AOI22_X1 i_3_43_128 (.A1(\buffer[11][4][3] [12]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][3] [12]), .ZN(n_3_43_115));
   AOI22_X1 i_3_43_129 (.A1(\buffer[13][4][3] [12]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][3] [12]), .ZN(n_3_43_116));
   NAND4_X1 i_3_43_130 (.A1(n_3_43_125), .A2(n_3_43_123), .A3(n_3_43_121), 
      .A4(n_3_43_117), .ZN(\output_filter[4][3] [13]));
   AOI221_X1 i_3_43_131 (.A(n_3_43_118), .B1(n_25), .B2(\buffer[0][4][3] [13]), 
      .C1(\buffer[12][4][3] [13]), .C2(n_27), .ZN(n_3_43_117));
   NAND4_X1 i_3_43_132 (.A1(n_3_43_124), .A2(n_3_43_122), .A3(n_3_43_120), 
      .A4(n_3_43_119), .ZN(n_3_43_118));
   AOI22_X1 i_3_43_133 (.A1(\buffer[15][4][3] [13]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][3] [13]), .ZN(n_3_43_119));
   AOI22_X1 i_3_43_134 (.A1(\buffer[10][4][3] [13]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][3] [13]), .ZN(n_3_43_120));
   AOI22_X1 i_3_43_135 (.A1(\buffer[6][4][3] [13]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][4][3] [13]), .ZN(n_3_43_121));
   AOI22_X1 i_3_43_136 (.A1(\buffer[9][4][3] [13]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][4][3] [13]), .ZN(n_3_43_122));
   AOI22_X1 i_3_43_137 (.A1(\buffer[14][4][3] [13]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][3] [13]), .ZN(n_3_43_123));
   AOI22_X1 i_3_43_138 (.A1(\buffer[11][4][3] [13]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][3] [13]), .ZN(n_3_43_124));
   AOI22_X1 i_3_43_139 (.A1(\buffer[13][4][3] [13]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][4][3] [13]), .ZN(n_3_43_125));
   NAND4_X1 i_3_43_140 (.A1(n_3_43_134), .A2(n_3_43_132), .A3(n_3_43_130), 
      .A4(n_3_43_126), .ZN(\output_filter[4][3] [14]));
   AOI221_X1 i_3_43_141 (.A(n_3_43_127), .B1(n_25), .B2(\buffer[0][4][3] [14]), 
      .C1(\buffer[12][4][3] [14]), .C2(n_27), .ZN(n_3_43_126));
   NAND4_X1 i_3_43_142 (.A1(n_3_43_133), .A2(n_3_43_131), .A3(n_3_43_129), 
      .A4(n_3_43_128), .ZN(n_3_43_127));
   AOI22_X1 i_3_43_143 (.A1(\buffer[15][4][3] [14]), .A2(n_22), .B1(n_16), 
      .B2(\buffer[8][4][3] [14]), .ZN(n_3_43_128));
   AOI22_X1 i_3_43_144 (.A1(\buffer[10][4][3] [14]), .A2(n_21), .B1(n_29), 
      .B2(\buffer[7][4][3] [14]), .ZN(n_3_43_129));
   AOI22_X1 i_3_43_145 (.A1(\buffer[6][4][3] [14]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][4][3] [14]), .ZN(n_3_43_130));
   AOI22_X1 i_3_43_146 (.A1(\buffer[9][4][3] [14]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][4][3] [14]), .ZN(n_3_43_131));
   AOI22_X1 i_3_43_147 (.A1(\buffer[14][4][3] [14]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][3] [14]), .ZN(n_3_43_132));
   AOI22_X1 i_3_43_148 (.A1(\buffer[11][4][3] [14]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][3] [14]), .ZN(n_3_43_133));
   AOI22_X1 i_3_43_149 (.A1(\buffer[13][4][3] [14]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][3] [14]), .ZN(n_3_43_134));
   NAND2_X1 i_3_43_150 (.A1(n_3_43_137), .A2(n_3_43_135), .ZN(
      \output_filter[4][3] [15]));
   AOI221_X1 i_3_43_151 (.A(n_3_43_136), .B1(n_31), .B2(\buffer[3][4][3] [15]), 
      .C1(\buffer[14][4][3] [15]), .C2(n_19), .ZN(n_3_43_135));
   NAND3_X1 i_3_43_152 (.A1(n_3_43_143), .A2(n_3_43_141), .A3(n_3_43_139), 
      .ZN(n_3_43_136));
   AOI221_X1 i_3_43_153 (.A(n_3_43_138), .B1(n_16), .B2(\buffer[8][4][3] [15]), 
      .C1(\buffer[13][4][3] [15]), .C2(n_26), .ZN(n_3_43_137));
   NAND3_X1 i_3_43_154 (.A1(n_3_43_144), .A2(n_3_43_142), .A3(n_3_43_140), 
      .ZN(n_3_43_138));
   AOI22_X1 i_3_43_155 (.A1(\buffer[11][4][3] [15]), .A2(n_17), .B1(n_24), 
      .B2(\buffer[2][4][3] [15]), .ZN(n_3_43_139));
   AOI22_X1 i_3_43_156 (.A1(\buffer[10][4][3] [15]), .A2(n_21), .B1(n_23), 
      .B2(\buffer[1][4][3] [15]), .ZN(n_3_43_140));
   AOI22_X1 i_3_43_157 (.A1(\buffer[6][4][3] [15]), .A2(n_28), .B1(n_18), 
      .B2(\buffer[5][4][3] [15]), .ZN(n_3_43_141));
   AOI22_X1 i_3_43_158 (.A1(\buffer[9][4][3] [15]), .A2(n_20), .B1(n_30), 
      .B2(\buffer[4][4][3] [15]), .ZN(n_3_43_142));
   AOI22_X1 i_3_43_159 (.A1(\buffer[7][4][3] [15]), .A2(n_29), .B1(n_25), 
      .B2(\buffer[0][4][3] [15]), .ZN(n_3_43_143));
   AOI22_X1 i_3_43_160 (.A1(\buffer[15][4][3] [15]), .A2(n_22), .B1(n_27), 
      .B2(\buffer[12][4][3] [15]), .ZN(n_3_43_144));
   NAND4_X1 i_4_42_0 (.A1(n_4_42_8), .A2(n_4_42_6), .A3(n_4_42_4), .A4(n_4_42_0), 
      .ZN(\output_filter[4][2] [0]));
   AOI221_X1 i_4_42_1 (.A(n_4_42_1), .B1(n_25), .B2(\buffer[0][4][2] [0]), 
      .C1(\buffer[12][4][2] [0]), .C2(n_27), .ZN(n_4_42_0));
   NAND4_X1 i_4_42_2 (.A1(n_4_42_7), .A2(n_4_42_5), .A3(n_4_42_3), .A4(n_4_42_2), 
      .ZN(n_4_42_1));
   AOI22_X1 i_4_42_3 (.A1(\buffer[15][4][2] [0]), .A2(n_22), .B1(n_29), .B2(
      \buffer[7][4][2] [0]), .ZN(n_4_42_2));
   AOI22_X1 i_4_42_4 (.A1(\buffer[10][4][2] [0]), .A2(n_21), .B1(n_16), .B2(
      \buffer[8][4][2] [0]), .ZN(n_4_42_3));
   AOI22_X1 i_4_42_5 (.A1(\buffer[6][4][2] [0]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][2] [0]), .ZN(n_4_42_4));
   AOI22_X1 i_4_42_6 (.A1(\buffer[9][4][2] [0]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][2] [0]), .ZN(n_4_42_5));
   AOI22_X1 i_4_42_7 (.A1(\buffer[14][4][2] [0]), .A2(n_19), .B1(n_23), .B2(
      \buffer[1][4][2] [0]), .ZN(n_4_42_6));
   AOI22_X1 i_4_42_8 (.A1(\buffer[11][4][2] [0]), .A2(n_17), .B1(n_18), .B2(
      \buffer[5][4][2] [0]), .ZN(n_4_42_7));
   AOI22_X1 i_4_42_9 (.A1(\buffer[13][4][2] [0]), .A2(n_26), .B1(n_24), .B2(
      \buffer[2][4][2] [0]), .ZN(n_4_42_8));
   NAND4_X1 i_4_42_10 (.A1(n_4_42_17), .A2(n_4_42_15), .A3(n_4_42_13), .A4(
      n_4_42_9), .ZN(\output_filter[4][2] [1]));
   AOI221_X1 i_4_42_11 (.A(n_4_42_10), .B1(n_25), .B2(\buffer[0][4][2] [1]), 
      .C1(\buffer[12][4][2] [1]), .C2(n_27), .ZN(n_4_42_9));
   NAND4_X1 i_4_42_12 (.A1(n_4_42_16), .A2(n_4_42_14), .A3(n_4_42_12), .A4(
      n_4_42_11), .ZN(n_4_42_10));
   AOI22_X1 i_4_42_13 (.A1(\buffer[15][4][2] [1]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][2] [1]), .ZN(n_4_42_11));
   AOI22_X1 i_4_42_14 (.A1(\buffer[10][4][2] [1]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][2] [1]), .ZN(n_4_42_12));
   AOI22_X1 i_4_42_15 (.A1(\buffer[6][4][2] [1]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][2] [1]), .ZN(n_4_42_13));
   AOI22_X1 i_4_42_16 (.A1(\buffer[9][4][2] [1]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][2] [1]), .ZN(n_4_42_14));
   AOI22_X1 i_4_42_17 (.A1(\buffer[14][4][2] [1]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][2] [1]), .ZN(n_4_42_15));
   AOI22_X1 i_4_42_18 (.A1(\buffer[11][4][2] [1]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][2] [1]), .ZN(n_4_42_16));
   AOI22_X1 i_4_42_19 (.A1(\buffer[13][4][2] [1]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][2] [1]), .ZN(n_4_42_17));
   NAND4_X1 i_4_42_20 (.A1(n_4_42_26), .A2(n_4_42_24), .A3(n_4_42_22), .A4(
      n_4_42_18), .ZN(\output_filter[4][2] [2]));
   AOI221_X1 i_4_42_21 (.A(n_4_42_19), .B1(n_25), .B2(\buffer[0][4][2] [2]), 
      .C1(\buffer[12][4][2] [2]), .C2(n_27), .ZN(n_4_42_18));
   NAND4_X1 i_4_42_22 (.A1(n_4_42_25), .A2(n_4_42_23), .A3(n_4_42_21), .A4(
      n_4_42_20), .ZN(n_4_42_19));
   AOI22_X1 i_4_42_23 (.A1(\buffer[15][4][2] [2]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][2] [2]), .ZN(n_4_42_20));
   AOI22_X1 i_4_42_24 (.A1(\buffer[10][4][2] [2]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][2] [2]), .ZN(n_4_42_21));
   AOI22_X1 i_4_42_25 (.A1(\buffer[6][4][2] [2]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][2] [2]), .ZN(n_4_42_22));
   AOI22_X1 i_4_42_26 (.A1(\buffer[9][4][2] [2]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][2] [2]), .ZN(n_4_42_23));
   AOI22_X1 i_4_42_27 (.A1(\buffer[14][4][2] [2]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][2] [2]), .ZN(n_4_42_24));
   AOI22_X1 i_4_42_28 (.A1(\buffer[11][4][2] [2]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][2] [2]), .ZN(n_4_42_25));
   AOI22_X1 i_4_42_29 (.A1(\buffer[13][4][2] [2]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][2] [2]), .ZN(n_4_42_26));
   NAND4_X1 i_4_42_30 (.A1(n_4_42_35), .A2(n_4_42_33), .A3(n_4_42_31), .A4(
      n_4_42_27), .ZN(\output_filter[4][2] [3]));
   AOI221_X1 i_4_42_31 (.A(n_4_42_28), .B1(n_25), .B2(\buffer[0][4][2] [3]), 
      .C1(\buffer[12][4][2] [3]), .C2(n_27), .ZN(n_4_42_27));
   NAND4_X1 i_4_42_32 (.A1(n_4_42_34), .A2(n_4_42_32), .A3(n_4_42_30), .A4(
      n_4_42_29), .ZN(n_4_42_28));
   AOI22_X1 i_4_42_33 (.A1(\buffer[15][4][2] [3]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][2] [3]), .ZN(n_4_42_29));
   AOI22_X1 i_4_42_34 (.A1(\buffer[10][4][2] [3]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][2] [3]), .ZN(n_4_42_30));
   AOI22_X1 i_4_42_35 (.A1(\buffer[6][4][2] [3]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][2] [3]), .ZN(n_4_42_31));
   AOI22_X1 i_4_42_36 (.A1(\buffer[9][4][2] [3]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][2] [3]), .ZN(n_4_42_32));
   AOI22_X1 i_4_42_37 (.A1(\buffer[14][4][2] [3]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][2] [3]), .ZN(n_4_42_33));
   AOI22_X1 i_4_42_38 (.A1(\buffer[11][4][2] [3]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][2] [3]), .ZN(n_4_42_34));
   AOI22_X1 i_4_42_39 (.A1(\buffer[13][4][2] [3]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][2] [3]), .ZN(n_4_42_35));
   NAND4_X1 i_4_42_40 (.A1(n_4_42_44), .A2(n_4_42_42), .A3(n_4_42_40), .A4(
      n_4_42_36), .ZN(\output_filter[4][2] [4]));
   AOI221_X1 i_4_42_41 (.A(n_4_42_37), .B1(n_25), .B2(\buffer[0][4][2] [4]), 
      .C1(\buffer[12][4][2] [4]), .C2(n_27), .ZN(n_4_42_36));
   NAND4_X1 i_4_42_42 (.A1(n_4_42_43), .A2(n_4_42_41), .A3(n_4_42_39), .A4(
      n_4_42_38), .ZN(n_4_42_37));
   AOI22_X1 i_4_42_43 (.A1(\buffer[15][4][2] [4]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][2] [4]), .ZN(n_4_42_38));
   AOI22_X1 i_4_42_44 (.A1(\buffer[10][4][2] [4]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][2] [4]), .ZN(n_4_42_39));
   AOI22_X1 i_4_42_45 (.A1(\buffer[6][4][2] [4]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][2] [4]), .ZN(n_4_42_40));
   AOI22_X1 i_4_42_46 (.A1(\buffer[9][4][2] [4]), .A2(n_20), .B1(n_24), .B2(
      \buffer[2][4][2] [4]), .ZN(n_4_42_41));
   AOI22_X1 i_4_42_47 (.A1(\buffer[14][4][2] [4]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][2] [4]), .ZN(n_4_42_42));
   AOI22_X1 i_4_42_48 (.A1(\buffer[11][4][2] [4]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][2] [4]), .ZN(n_4_42_43));
   AOI22_X1 i_4_42_49 (.A1(\buffer[13][4][2] [4]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][4][2] [4]), .ZN(n_4_42_44));
   NAND4_X1 i_4_42_50 (.A1(n_4_42_53), .A2(n_4_42_51), .A3(n_4_42_49), .A4(
      n_4_42_45), .ZN(\output_filter[4][2] [5]));
   AOI221_X1 i_4_42_51 (.A(n_4_42_46), .B1(n_25), .B2(\buffer[0][4][2] [5]), 
      .C1(\buffer[12][4][2] [5]), .C2(n_27), .ZN(n_4_42_45));
   NAND4_X1 i_4_42_52 (.A1(n_4_42_52), .A2(n_4_42_50), .A3(n_4_42_48), .A4(
      n_4_42_47), .ZN(n_4_42_46));
   AOI22_X1 i_4_42_53 (.A1(\buffer[15][4][2] [5]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][2] [5]), .ZN(n_4_42_47));
   AOI22_X1 i_4_42_54 (.A1(\buffer[10][4][2] [5]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][2] [5]), .ZN(n_4_42_48));
   AOI22_X1 i_4_42_55 (.A1(\buffer[6][4][2] [5]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][2] [5]), .ZN(n_4_42_49));
   AOI22_X1 i_4_42_56 (.A1(\buffer[9][4][2] [5]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][2] [5]), .ZN(n_4_42_50));
   AOI22_X1 i_4_42_57 (.A1(\buffer[14][4][2] [5]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][2] [5]), .ZN(n_4_42_51));
   AOI22_X1 i_4_42_58 (.A1(\buffer[11][4][2] [5]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][2] [5]), .ZN(n_4_42_52));
   AOI22_X1 i_4_42_59 (.A1(\buffer[13][4][2] [5]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][2] [5]), .ZN(n_4_42_53));
   NAND4_X1 i_4_42_60 (.A1(n_4_42_62), .A2(n_4_42_60), .A3(n_4_42_58), .A4(
      n_4_42_54), .ZN(\output_filter[4][2] [6]));
   AOI221_X1 i_4_42_61 (.A(n_4_42_55), .B1(n_25), .B2(\buffer[0][4][2] [6]), 
      .C1(\buffer[12][4][2] [6]), .C2(n_27), .ZN(n_4_42_54));
   NAND4_X1 i_4_42_62 (.A1(n_4_42_61), .A2(n_4_42_59), .A3(n_4_42_57), .A4(
      n_4_42_56), .ZN(n_4_42_55));
   AOI22_X1 i_4_42_63 (.A1(\buffer[15][4][2] [6]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][2] [6]), .ZN(n_4_42_56));
   AOI22_X1 i_4_42_64 (.A1(\buffer[10][4][2] [6]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][2] [6]), .ZN(n_4_42_57));
   AOI22_X1 i_4_42_65 (.A1(\buffer[6][4][2] [6]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][2] [6]), .ZN(n_4_42_58));
   AOI22_X1 i_4_42_66 (.A1(\buffer[9][4][2] [6]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][2] [6]), .ZN(n_4_42_59));
   AOI22_X1 i_4_42_67 (.A1(\buffer[14][4][2] [6]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][2] [6]), .ZN(n_4_42_60));
   AOI22_X1 i_4_42_68 (.A1(\buffer[11][4][2] [6]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][2] [6]), .ZN(n_4_42_61));
   AOI22_X1 i_4_42_69 (.A1(\buffer[13][4][2] [6]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][2] [6]), .ZN(n_4_42_62));
   NAND4_X1 i_4_42_70 (.A1(n_4_42_71), .A2(n_4_42_69), .A3(n_4_42_67), .A4(
      n_4_42_63), .ZN(\output_filter[4][2] [7]));
   AOI221_X1 i_4_42_71 (.A(n_4_42_64), .B1(n_25), .B2(\buffer[0][4][2] [7]), 
      .C1(\buffer[12][4][2] [7]), .C2(n_27), .ZN(n_4_42_63));
   NAND4_X1 i_4_42_72 (.A1(n_4_42_70), .A2(n_4_42_68), .A3(n_4_42_66), .A4(
      n_4_42_65), .ZN(n_4_42_64));
   AOI22_X1 i_4_42_73 (.A1(\buffer[15][4][2] [7]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][2] [7]), .ZN(n_4_42_65));
   AOI22_X1 i_4_42_74 (.A1(\buffer[10][4][2] [7]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][2] [7]), .ZN(n_4_42_66));
   AOI22_X1 i_4_42_75 (.A1(\buffer[6][4][2] [7]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][2] [7]), .ZN(n_4_42_67));
   AOI22_X1 i_4_42_76 (.A1(\buffer[9][4][2] [7]), .A2(n_20), .B1(n_24), .B2(
      \buffer[2][4][2] [7]), .ZN(n_4_42_68));
   AOI22_X1 i_4_42_77 (.A1(\buffer[14][4][2] [7]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][2] [7]), .ZN(n_4_42_69));
   AOI22_X1 i_4_42_78 (.A1(\buffer[11][4][2] [7]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][2] [7]), .ZN(n_4_42_70));
   AOI22_X1 i_4_42_79 (.A1(\buffer[13][4][2] [7]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][4][2] [7]), .ZN(n_4_42_71));
   NAND4_X1 i_4_42_80 (.A1(n_4_42_80), .A2(n_4_42_78), .A3(n_4_42_76), .A4(
      n_4_42_72), .ZN(\output_filter[4][2] [8]));
   AOI221_X1 i_4_42_81 (.A(n_4_42_73), .B1(n_25), .B2(\buffer[0][4][2] [8]), 
      .C1(\buffer[12][4][2] [8]), .C2(n_27), .ZN(n_4_42_72));
   NAND4_X1 i_4_42_82 (.A1(n_4_42_79), .A2(n_4_42_77), .A3(n_4_42_75), .A4(
      n_4_42_74), .ZN(n_4_42_73));
   AOI22_X1 i_4_42_83 (.A1(\buffer[15][4][2] [8]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][2] [8]), .ZN(n_4_42_74));
   AOI22_X1 i_4_42_84 (.A1(\buffer[10][4][2] [8]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][2] [8]), .ZN(n_4_42_75));
   AOI22_X1 i_4_42_85 (.A1(\buffer[6][4][2] [8]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][2] [8]), .ZN(n_4_42_76));
   AOI22_X1 i_4_42_86 (.A1(\buffer[9][4][2] [8]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][2] [8]), .ZN(n_4_42_77));
   AOI22_X1 i_4_42_87 (.A1(\buffer[14][4][2] [8]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][2] [8]), .ZN(n_4_42_78));
   AOI22_X1 i_4_42_88 (.A1(\buffer[11][4][2] [8]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][2] [8]), .ZN(n_4_42_79));
   AOI22_X1 i_4_42_89 (.A1(\buffer[13][4][2] [8]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][2] [8]), .ZN(n_4_42_80));
   NAND4_X1 i_4_42_90 (.A1(n_4_42_89), .A2(n_4_42_87), .A3(n_4_42_85), .A4(
      n_4_42_81), .ZN(\output_filter[4][2] [9]));
   AOI221_X1 i_4_42_91 (.A(n_4_42_82), .B1(n_25), .B2(\buffer[0][4][2] [9]), 
      .C1(\buffer[12][4][2] [9]), .C2(n_27), .ZN(n_4_42_81));
   NAND4_X1 i_4_42_92 (.A1(n_4_42_88), .A2(n_4_42_86), .A3(n_4_42_84), .A4(
      n_4_42_83), .ZN(n_4_42_82));
   AOI22_X1 i_4_42_93 (.A1(\buffer[15][4][2] [9]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][2] [9]), .ZN(n_4_42_83));
   AOI22_X1 i_4_42_94 (.A1(\buffer[10][4][2] [9]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][2] [9]), .ZN(n_4_42_84));
   AOI22_X1 i_4_42_95 (.A1(\buffer[6][4][2] [9]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][2] [9]), .ZN(n_4_42_85));
   AOI22_X1 i_4_42_96 (.A1(\buffer[9][4][2] [9]), .A2(n_20), .B1(n_24), .B2(
      \buffer[2][4][2] [9]), .ZN(n_4_42_86));
   AOI22_X1 i_4_42_97 (.A1(\buffer[14][4][2] [9]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][2] [9]), .ZN(n_4_42_87));
   AOI22_X1 i_4_42_98 (.A1(\buffer[11][4][2] [9]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][2] [9]), .ZN(n_4_42_88));
   AOI22_X1 i_4_42_99 (.A1(\buffer[13][4][2] [9]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][4][2] [9]), .ZN(n_4_42_89));
   NAND4_X1 i_4_42_100 (.A1(n_4_42_98), .A2(n_4_42_96), .A3(n_4_42_94), .A4(
      n_4_42_90), .ZN(\output_filter[4][2] [10]));
   AOI221_X1 i_4_42_101 (.A(n_4_42_91), .B1(n_25), .B2(\buffer[0][4][2] [10]), 
      .C1(\buffer[12][4][2] [10]), .C2(n_27), .ZN(n_4_42_90));
   NAND4_X1 i_4_42_102 (.A1(n_4_42_97), .A2(n_4_42_95), .A3(n_4_42_93), .A4(
      n_4_42_92), .ZN(n_4_42_91));
   AOI22_X1 i_4_42_103 (.A1(\buffer[15][4][2] [10]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][2] [10]), .ZN(n_4_42_92));
   AOI22_X1 i_4_42_104 (.A1(\buffer[10][4][2] [10]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][2] [10]), .ZN(n_4_42_93));
   AOI22_X1 i_4_42_105 (.A1(\buffer[6][4][2] [10]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][4][2] [10]), .ZN(n_4_42_94));
   AOI22_X1 i_4_42_106 (.A1(\buffer[9][4][2] [10]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][4][2] [10]), .ZN(n_4_42_95));
   AOI22_X1 i_4_42_107 (.A1(\buffer[14][4][2] [10]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][2] [10]), .ZN(n_4_42_96));
   AOI22_X1 i_4_42_108 (.A1(\buffer[11][4][2] [10]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][2] [10]), .ZN(n_4_42_97));
   AOI22_X1 i_4_42_109 (.A1(\buffer[13][4][2] [10]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][2] [10]), .ZN(n_4_42_98));
   NAND4_X1 i_4_42_110 (.A1(n_4_42_107), .A2(n_4_42_105), .A3(n_4_42_103), 
      .A4(n_4_42_99), .ZN(\output_filter[4][2] [11]));
   AOI221_X1 i_4_42_111 (.A(n_4_42_100), .B1(n_25), .B2(\buffer[0][4][2] [11]), 
      .C1(\buffer[12][4][2] [11]), .C2(n_27), .ZN(n_4_42_99));
   NAND4_X1 i_4_42_112 (.A1(n_4_42_106), .A2(n_4_42_104), .A3(n_4_42_102), 
      .A4(n_4_42_101), .ZN(n_4_42_100));
   AOI22_X1 i_4_42_113 (.A1(\buffer[15][4][2] [11]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][2] [11]), .ZN(n_4_42_101));
   AOI22_X1 i_4_42_114 (.A1(\buffer[10][4][2] [11]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][2] [11]), .ZN(n_4_42_102));
   AOI22_X1 i_4_42_115 (.A1(\buffer[6][4][2] [11]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][4][2] [11]), .ZN(n_4_42_103));
   AOI22_X1 i_4_42_116 (.A1(\buffer[9][4][2] [11]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][4][2] [11]), .ZN(n_4_42_104));
   AOI22_X1 i_4_42_117 (.A1(\buffer[14][4][2] [11]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][2] [11]), .ZN(n_4_42_105));
   AOI22_X1 i_4_42_118 (.A1(\buffer[11][4][2] [11]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][2] [11]), .ZN(n_4_42_106));
   AOI22_X1 i_4_42_119 (.A1(\buffer[13][4][2] [11]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][4][2] [11]), .ZN(n_4_42_107));
   NAND4_X1 i_4_42_120 (.A1(n_4_42_116), .A2(n_4_42_114), .A3(n_4_42_112), 
      .A4(n_4_42_108), .ZN(\output_filter[4][2] [12]));
   AOI221_X1 i_4_42_121 (.A(n_4_42_109), .B1(n_25), .B2(\buffer[0][4][2] [12]), 
      .C1(\buffer[12][4][2] [12]), .C2(n_27), .ZN(n_4_42_108));
   NAND4_X1 i_4_42_122 (.A1(n_4_42_115), .A2(n_4_42_113), .A3(n_4_42_111), 
      .A4(n_4_42_110), .ZN(n_4_42_109));
   AOI22_X1 i_4_42_123 (.A1(\buffer[15][4][2] [12]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][2] [12]), .ZN(n_4_42_110));
   AOI22_X1 i_4_42_124 (.A1(\buffer[10][4][2] [12]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][2] [12]), .ZN(n_4_42_111));
   AOI22_X1 i_4_42_125 (.A1(\buffer[6][4][2] [12]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][4][2] [12]), .ZN(n_4_42_112));
   AOI22_X1 i_4_42_126 (.A1(\buffer[9][4][2] [12]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][4][2] [12]), .ZN(n_4_42_113));
   AOI22_X1 i_4_42_127 (.A1(\buffer[14][4][2] [12]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][2] [12]), .ZN(n_4_42_114));
   AOI22_X1 i_4_42_128 (.A1(\buffer[11][4][2] [12]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][2] [12]), .ZN(n_4_42_115));
   AOI22_X1 i_4_42_129 (.A1(\buffer[13][4][2] [12]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][2] [12]), .ZN(n_4_42_116));
   NAND4_X1 i_4_42_130 (.A1(n_4_42_125), .A2(n_4_42_123), .A3(n_4_42_121), 
      .A4(n_4_42_117), .ZN(\output_filter[4][2] [13]));
   AOI221_X1 i_4_42_131 (.A(n_4_42_118), .B1(n_25), .B2(\buffer[0][4][2] [13]), 
      .C1(\buffer[12][4][2] [13]), .C2(n_27), .ZN(n_4_42_117));
   NAND4_X1 i_4_42_132 (.A1(n_4_42_124), .A2(n_4_42_122), .A3(n_4_42_120), 
      .A4(n_4_42_119), .ZN(n_4_42_118));
   AOI22_X1 i_4_42_133 (.A1(\buffer[15][4][2] [13]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][2] [13]), .ZN(n_4_42_119));
   AOI22_X1 i_4_42_134 (.A1(\buffer[10][4][2] [13]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][2] [13]), .ZN(n_4_42_120));
   AOI22_X1 i_4_42_135 (.A1(\buffer[6][4][2] [13]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][4][2] [13]), .ZN(n_4_42_121));
   AOI22_X1 i_4_42_136 (.A1(\buffer[9][4][2] [13]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][4][2] [13]), .ZN(n_4_42_122));
   AOI22_X1 i_4_42_137 (.A1(\buffer[14][4][2] [13]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][2] [13]), .ZN(n_4_42_123));
   AOI22_X1 i_4_42_138 (.A1(\buffer[11][4][2] [13]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][2] [13]), .ZN(n_4_42_124));
   AOI22_X1 i_4_42_139 (.A1(\buffer[13][4][2] [13]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][4][2] [13]), .ZN(n_4_42_125));
   NAND4_X1 i_4_42_140 (.A1(n_4_42_134), .A2(n_4_42_132), .A3(n_4_42_130), 
      .A4(n_4_42_126), .ZN(\output_filter[4][2] [14]));
   AOI221_X1 i_4_42_141 (.A(n_4_42_127), .B1(n_25), .B2(\buffer[0][4][2] [14]), 
      .C1(\buffer[12][4][2] [14]), .C2(n_27), .ZN(n_4_42_126));
   NAND4_X1 i_4_42_142 (.A1(n_4_42_133), .A2(n_4_42_131), .A3(n_4_42_129), 
      .A4(n_4_42_128), .ZN(n_4_42_127));
   AOI22_X1 i_4_42_143 (.A1(\buffer[15][4][2] [14]), .A2(n_22), .B1(n_16), 
      .B2(\buffer[8][4][2] [14]), .ZN(n_4_42_128));
   AOI22_X1 i_4_42_144 (.A1(\buffer[10][4][2] [14]), .A2(n_21), .B1(n_29), 
      .B2(\buffer[7][4][2] [14]), .ZN(n_4_42_129));
   AOI22_X1 i_4_42_145 (.A1(\buffer[6][4][2] [14]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][4][2] [14]), .ZN(n_4_42_130));
   AOI22_X1 i_4_42_146 (.A1(\buffer[9][4][2] [14]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][4][2] [14]), .ZN(n_4_42_131));
   AOI22_X1 i_4_42_147 (.A1(\buffer[14][4][2] [14]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][2] [14]), .ZN(n_4_42_132));
   AOI22_X1 i_4_42_148 (.A1(\buffer[11][4][2] [14]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][2] [14]), .ZN(n_4_42_133));
   AOI22_X1 i_4_42_149 (.A1(\buffer[13][4][2] [14]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][2] [14]), .ZN(n_4_42_134));
   NAND2_X1 i_4_42_150 (.A1(n_4_42_137), .A2(n_4_42_135), .ZN(
      \output_filter[4][2] [15]));
   AOI221_X1 i_4_42_151 (.A(n_4_42_136), .B1(n_31), .B2(\buffer[3][4][2] [15]), 
      .C1(\buffer[14][4][2] [15]), .C2(n_19), .ZN(n_4_42_135));
   NAND3_X1 i_4_42_152 (.A1(n_4_42_143), .A2(n_4_42_141), .A3(n_4_42_139), 
      .ZN(n_4_42_136));
   AOI221_X1 i_4_42_153 (.A(n_4_42_138), .B1(n_16), .B2(\buffer[8][4][2] [15]), 
      .C1(\buffer[13][4][2] [15]), .C2(n_26), .ZN(n_4_42_137));
   NAND3_X1 i_4_42_154 (.A1(n_4_42_144), .A2(n_4_42_142), .A3(n_4_42_140), 
      .ZN(n_4_42_138));
   AOI22_X1 i_4_42_155 (.A1(\buffer[11][4][2] [15]), .A2(n_17), .B1(n_24), 
      .B2(\buffer[2][4][2] [15]), .ZN(n_4_42_139));
   AOI22_X1 i_4_42_156 (.A1(\buffer[10][4][2] [15]), .A2(n_21), .B1(n_23), 
      .B2(\buffer[1][4][2] [15]), .ZN(n_4_42_140));
   AOI22_X1 i_4_42_157 (.A1(\buffer[6][4][2] [15]), .A2(n_28), .B1(n_18), 
      .B2(\buffer[5][4][2] [15]), .ZN(n_4_42_141));
   AOI22_X1 i_4_42_158 (.A1(\buffer[9][4][2] [15]), .A2(n_20), .B1(n_30), 
      .B2(\buffer[4][4][2] [15]), .ZN(n_4_42_142));
   AOI22_X1 i_4_42_159 (.A1(\buffer[7][4][2] [15]), .A2(n_29), .B1(n_25), 
      .B2(\buffer[0][4][2] [15]), .ZN(n_4_42_143));
   AOI22_X1 i_4_42_160 (.A1(\buffer[15][4][2] [15]), .A2(n_22), .B1(n_27), 
      .B2(\buffer[12][4][2] [15]), .ZN(n_4_42_144));
   NAND4_X1 i_5_41_0 (.A1(n_5_41_8), .A2(n_5_41_6), .A3(n_5_41_4), .A4(n_5_41_0), 
      .ZN(\output_filter[4][1] [0]));
   AOI221_X1 i_5_41_1 (.A(n_5_41_1), .B1(n_25), .B2(\buffer[0][4][1] [0]), 
      .C1(\buffer[12][4][1] [0]), .C2(n_27), .ZN(n_5_41_0));
   NAND4_X1 i_5_41_2 (.A1(n_5_41_7), .A2(n_5_41_5), .A3(n_5_41_3), .A4(n_5_41_2), 
      .ZN(n_5_41_1));
   AOI22_X1 i_5_41_3 (.A1(\buffer[15][4][1] [0]), .A2(n_22), .B1(n_29), .B2(
      \buffer[7][4][1] [0]), .ZN(n_5_41_2));
   AOI22_X1 i_5_41_4 (.A1(\buffer[10][4][1] [0]), .A2(n_21), .B1(n_16), .B2(
      \buffer[8][4][1] [0]), .ZN(n_5_41_3));
   AOI22_X1 i_5_41_5 (.A1(\buffer[6][4][1] [0]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][1] [0]), .ZN(n_5_41_4));
   AOI22_X1 i_5_41_6 (.A1(\buffer[9][4][1] [0]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][1] [0]), .ZN(n_5_41_5));
   AOI22_X1 i_5_41_7 (.A1(\buffer[14][4][1] [0]), .A2(n_19), .B1(n_23), .B2(
      \buffer[1][4][1] [0]), .ZN(n_5_41_6));
   AOI22_X1 i_5_41_8 (.A1(\buffer[11][4][1] [0]), .A2(n_17), .B1(n_18), .B2(
      \buffer[5][4][1] [0]), .ZN(n_5_41_7));
   AOI22_X1 i_5_41_9 (.A1(\buffer[13][4][1] [0]), .A2(n_26), .B1(n_24), .B2(
      \buffer[2][4][1] [0]), .ZN(n_5_41_8));
   NAND4_X1 i_5_41_10 (.A1(n_5_41_17), .A2(n_5_41_15), .A3(n_5_41_13), .A4(
      n_5_41_9), .ZN(\output_filter[4][1] [1]));
   AOI221_X1 i_5_41_11 (.A(n_5_41_10), .B1(n_25), .B2(\buffer[0][4][1] [1]), 
      .C1(\buffer[12][4][1] [1]), .C2(n_27), .ZN(n_5_41_9));
   NAND4_X1 i_5_41_12 (.A1(n_5_41_16), .A2(n_5_41_14), .A3(n_5_41_12), .A4(
      n_5_41_11), .ZN(n_5_41_10));
   AOI22_X1 i_5_41_13 (.A1(\buffer[15][4][1] [1]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][1] [1]), .ZN(n_5_41_11));
   AOI22_X1 i_5_41_14 (.A1(\buffer[10][4][1] [1]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][1] [1]), .ZN(n_5_41_12));
   AOI22_X1 i_5_41_15 (.A1(\buffer[6][4][1] [1]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][1] [1]), .ZN(n_5_41_13));
   AOI22_X1 i_5_41_16 (.A1(\buffer[9][4][1] [1]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][1] [1]), .ZN(n_5_41_14));
   AOI22_X1 i_5_41_17 (.A1(\buffer[14][4][1] [1]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][1] [1]), .ZN(n_5_41_15));
   AOI22_X1 i_5_41_18 (.A1(\buffer[11][4][1] [1]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][1] [1]), .ZN(n_5_41_16));
   AOI22_X1 i_5_41_19 (.A1(\buffer[13][4][1] [1]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][1] [1]), .ZN(n_5_41_17));
   NAND4_X1 i_5_41_20 (.A1(n_5_41_26), .A2(n_5_41_24), .A3(n_5_41_22), .A4(
      n_5_41_18), .ZN(\output_filter[4][1] [2]));
   AOI221_X1 i_5_41_21 (.A(n_5_41_19), .B1(n_25), .B2(\buffer[0][4][1] [2]), 
      .C1(\buffer[12][4][1] [2]), .C2(n_27), .ZN(n_5_41_18));
   NAND4_X1 i_5_41_22 (.A1(n_5_41_25), .A2(n_5_41_23), .A3(n_5_41_21), .A4(
      n_5_41_20), .ZN(n_5_41_19));
   AOI22_X1 i_5_41_23 (.A1(\buffer[15][4][1] [2]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][1] [2]), .ZN(n_5_41_20));
   AOI22_X1 i_5_41_24 (.A1(\buffer[10][4][1] [2]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][1] [2]), .ZN(n_5_41_21));
   AOI22_X1 i_5_41_25 (.A1(\buffer[6][4][1] [2]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][1] [2]), .ZN(n_5_41_22));
   AOI22_X1 i_5_41_26 (.A1(\buffer[9][4][1] [2]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][1] [2]), .ZN(n_5_41_23));
   AOI22_X1 i_5_41_27 (.A1(\buffer[14][4][1] [2]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][1] [2]), .ZN(n_5_41_24));
   AOI22_X1 i_5_41_28 (.A1(\buffer[11][4][1] [2]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][1] [2]), .ZN(n_5_41_25));
   AOI22_X1 i_5_41_29 (.A1(\buffer[13][4][1] [2]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][1] [2]), .ZN(n_5_41_26));
   NAND4_X1 i_5_41_30 (.A1(n_5_41_35), .A2(n_5_41_33), .A3(n_5_41_31), .A4(
      n_5_41_27), .ZN(\output_filter[4][1] [3]));
   AOI221_X1 i_5_41_31 (.A(n_5_41_28), .B1(n_25), .B2(\buffer[0][4][1] [3]), 
      .C1(\buffer[12][4][1] [3]), .C2(n_27), .ZN(n_5_41_27));
   NAND4_X1 i_5_41_32 (.A1(n_5_41_34), .A2(n_5_41_32), .A3(n_5_41_30), .A4(
      n_5_41_29), .ZN(n_5_41_28));
   AOI22_X1 i_5_41_33 (.A1(\buffer[15][4][1] [3]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][1] [3]), .ZN(n_5_41_29));
   AOI22_X1 i_5_41_34 (.A1(\buffer[10][4][1] [3]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][1] [3]), .ZN(n_5_41_30));
   AOI22_X1 i_5_41_35 (.A1(\buffer[6][4][1] [3]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][1] [3]), .ZN(n_5_41_31));
   AOI22_X1 i_5_41_36 (.A1(\buffer[9][4][1] [3]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][1] [3]), .ZN(n_5_41_32));
   AOI22_X1 i_5_41_37 (.A1(\buffer[14][4][1] [3]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][1] [3]), .ZN(n_5_41_33));
   AOI22_X1 i_5_41_38 (.A1(\buffer[11][4][1] [3]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][1] [3]), .ZN(n_5_41_34));
   AOI22_X1 i_5_41_39 (.A1(\buffer[13][4][1] [3]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][1] [3]), .ZN(n_5_41_35));
   NAND4_X1 i_5_41_40 (.A1(n_5_41_44), .A2(n_5_41_42), .A3(n_5_41_40), .A4(
      n_5_41_36), .ZN(\output_filter[4][1] [4]));
   AOI221_X1 i_5_41_41 (.A(n_5_41_37), .B1(n_25), .B2(\buffer[0][4][1] [4]), 
      .C1(\buffer[12][4][1] [4]), .C2(n_27), .ZN(n_5_41_36));
   NAND4_X1 i_5_41_42 (.A1(n_5_41_43), .A2(n_5_41_41), .A3(n_5_41_39), .A4(
      n_5_41_38), .ZN(n_5_41_37));
   AOI22_X1 i_5_41_43 (.A1(\buffer[15][4][1] [4]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][1] [4]), .ZN(n_5_41_38));
   AOI22_X1 i_5_41_44 (.A1(\buffer[10][4][1] [4]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][1] [4]), .ZN(n_5_41_39));
   AOI22_X1 i_5_41_45 (.A1(\buffer[6][4][1] [4]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][1] [4]), .ZN(n_5_41_40));
   AOI22_X1 i_5_41_46 (.A1(\buffer[9][4][1] [4]), .A2(n_20), .B1(n_24), .B2(
      \buffer[2][4][1] [4]), .ZN(n_5_41_41));
   AOI22_X1 i_5_41_47 (.A1(\buffer[14][4][1] [4]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][1] [4]), .ZN(n_5_41_42));
   AOI22_X1 i_5_41_48 (.A1(\buffer[11][4][1] [4]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][1] [4]), .ZN(n_5_41_43));
   AOI22_X1 i_5_41_49 (.A1(\buffer[13][4][1] [4]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][4][1] [4]), .ZN(n_5_41_44));
   NAND4_X1 i_5_41_50 (.A1(n_5_41_53), .A2(n_5_41_51), .A3(n_5_41_49), .A4(
      n_5_41_45), .ZN(\output_filter[4][1] [5]));
   AOI221_X1 i_5_41_51 (.A(n_5_41_46), .B1(n_25), .B2(\buffer[0][4][1] [5]), 
      .C1(\buffer[12][4][1] [5]), .C2(n_27), .ZN(n_5_41_45));
   NAND4_X1 i_5_41_52 (.A1(n_5_41_52), .A2(n_5_41_50), .A3(n_5_41_48), .A4(
      n_5_41_47), .ZN(n_5_41_46));
   AOI22_X1 i_5_41_53 (.A1(\buffer[15][4][1] [5]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][1] [5]), .ZN(n_5_41_47));
   AOI22_X1 i_5_41_54 (.A1(\buffer[10][4][1] [5]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][1] [5]), .ZN(n_5_41_48));
   AOI22_X1 i_5_41_55 (.A1(\buffer[6][4][1] [5]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][1] [5]), .ZN(n_5_41_49));
   AOI22_X1 i_5_41_56 (.A1(\buffer[9][4][1] [5]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][1] [5]), .ZN(n_5_41_50));
   AOI22_X1 i_5_41_57 (.A1(\buffer[14][4][1] [5]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][1] [5]), .ZN(n_5_41_51));
   AOI22_X1 i_5_41_58 (.A1(\buffer[11][4][1] [5]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][1] [5]), .ZN(n_5_41_52));
   AOI22_X1 i_5_41_59 (.A1(\buffer[13][4][1] [5]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][1] [5]), .ZN(n_5_41_53));
   NAND4_X1 i_5_41_60 (.A1(n_5_41_62), .A2(n_5_41_60), .A3(n_5_41_58), .A4(
      n_5_41_54), .ZN(\output_filter[4][1] [6]));
   AOI221_X1 i_5_41_61 (.A(n_5_41_55), .B1(n_25), .B2(\buffer[0][4][1] [6]), 
      .C1(\buffer[12][4][1] [6]), .C2(n_27), .ZN(n_5_41_54));
   NAND4_X1 i_5_41_62 (.A1(n_5_41_61), .A2(n_5_41_59), .A3(n_5_41_57), .A4(
      n_5_41_56), .ZN(n_5_41_55));
   AOI22_X1 i_5_41_63 (.A1(\buffer[15][4][1] [6]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][1] [6]), .ZN(n_5_41_56));
   AOI22_X1 i_5_41_64 (.A1(\buffer[10][4][1] [6]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][1] [6]), .ZN(n_5_41_57));
   AOI22_X1 i_5_41_65 (.A1(\buffer[6][4][1] [6]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][1] [6]), .ZN(n_5_41_58));
   AOI22_X1 i_5_41_66 (.A1(\buffer[9][4][1] [6]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][1] [6]), .ZN(n_5_41_59));
   AOI22_X1 i_5_41_67 (.A1(\buffer[14][4][1] [6]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][1] [6]), .ZN(n_5_41_60));
   AOI22_X1 i_5_41_68 (.A1(\buffer[11][4][1] [6]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][1] [6]), .ZN(n_5_41_61));
   AOI22_X1 i_5_41_69 (.A1(\buffer[13][4][1] [6]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][1] [6]), .ZN(n_5_41_62));
   NAND4_X1 i_5_41_70 (.A1(n_5_41_71), .A2(n_5_41_69), .A3(n_5_41_67), .A4(
      n_5_41_63), .ZN(\output_filter[4][1] [7]));
   AOI221_X1 i_5_41_71 (.A(n_5_41_64), .B1(n_25), .B2(\buffer[0][4][1] [7]), 
      .C1(\buffer[12][4][1] [7]), .C2(n_27), .ZN(n_5_41_63));
   NAND4_X1 i_5_41_72 (.A1(n_5_41_70), .A2(n_5_41_68), .A3(n_5_41_66), .A4(
      n_5_41_65), .ZN(n_5_41_64));
   AOI22_X1 i_5_41_73 (.A1(\buffer[15][4][1] [7]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][1] [7]), .ZN(n_5_41_65));
   AOI22_X1 i_5_41_74 (.A1(\buffer[10][4][1] [7]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][1] [7]), .ZN(n_5_41_66));
   AOI22_X1 i_5_41_75 (.A1(\buffer[6][4][1] [7]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][1] [7]), .ZN(n_5_41_67));
   AOI22_X1 i_5_41_76 (.A1(\buffer[9][4][1] [7]), .A2(n_20), .B1(n_24), .B2(
      \buffer[2][4][1] [7]), .ZN(n_5_41_68));
   AOI22_X1 i_5_41_77 (.A1(\buffer[14][4][1] [7]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][1] [7]), .ZN(n_5_41_69));
   AOI22_X1 i_5_41_78 (.A1(\buffer[11][4][1] [7]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][1] [7]), .ZN(n_5_41_70));
   AOI22_X1 i_5_41_79 (.A1(\buffer[13][4][1] [7]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][4][1] [7]), .ZN(n_5_41_71));
   NAND4_X1 i_5_41_80 (.A1(n_5_41_80), .A2(n_5_41_78), .A3(n_5_41_76), .A4(
      n_5_41_72), .ZN(\output_filter[4][1] [8]));
   AOI221_X1 i_5_41_81 (.A(n_5_41_73), .B1(n_25), .B2(\buffer[0][4][1] [8]), 
      .C1(\buffer[12][4][1] [8]), .C2(n_27), .ZN(n_5_41_72));
   NAND4_X1 i_5_41_82 (.A1(n_5_41_79), .A2(n_5_41_77), .A3(n_5_41_75), .A4(
      n_5_41_74), .ZN(n_5_41_73));
   AOI22_X1 i_5_41_83 (.A1(\buffer[15][4][1] [8]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][1] [8]), .ZN(n_5_41_74));
   AOI22_X1 i_5_41_84 (.A1(\buffer[10][4][1] [8]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][1] [8]), .ZN(n_5_41_75));
   AOI22_X1 i_5_41_85 (.A1(\buffer[6][4][1] [8]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][1] [8]), .ZN(n_5_41_76));
   AOI22_X1 i_5_41_86 (.A1(\buffer[9][4][1] [8]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][1] [8]), .ZN(n_5_41_77));
   AOI22_X1 i_5_41_87 (.A1(\buffer[14][4][1] [8]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][1] [8]), .ZN(n_5_41_78));
   AOI22_X1 i_5_41_88 (.A1(\buffer[11][4][1] [8]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][1] [8]), .ZN(n_5_41_79));
   AOI22_X1 i_5_41_89 (.A1(\buffer[13][4][1] [8]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][1] [8]), .ZN(n_5_41_80));
   NAND4_X1 i_5_41_90 (.A1(n_5_41_89), .A2(n_5_41_87), .A3(n_5_41_85), .A4(
      n_5_41_81), .ZN(\output_filter[4][1] [9]));
   AOI221_X1 i_5_41_91 (.A(n_5_41_82), .B1(n_25), .B2(\buffer[0][4][1] [9]), 
      .C1(\buffer[12][4][1] [9]), .C2(n_27), .ZN(n_5_41_81));
   NAND4_X1 i_5_41_92 (.A1(n_5_41_88), .A2(n_5_41_86), .A3(n_5_41_84), .A4(
      n_5_41_83), .ZN(n_5_41_82));
   AOI22_X1 i_5_41_93 (.A1(\buffer[15][4][1] [9]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][1] [9]), .ZN(n_5_41_83));
   AOI22_X1 i_5_41_94 (.A1(\buffer[10][4][1] [9]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][1] [9]), .ZN(n_5_41_84));
   AOI22_X1 i_5_41_95 (.A1(\buffer[6][4][1] [9]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][1] [9]), .ZN(n_5_41_85));
   AOI22_X1 i_5_41_96 (.A1(\buffer[9][4][1] [9]), .A2(n_20), .B1(n_24), .B2(
      \buffer[2][4][1] [9]), .ZN(n_5_41_86));
   AOI22_X1 i_5_41_97 (.A1(\buffer[14][4][1] [9]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][1] [9]), .ZN(n_5_41_87));
   AOI22_X1 i_5_41_98 (.A1(\buffer[11][4][1] [9]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][1] [9]), .ZN(n_5_41_88));
   AOI22_X1 i_5_41_99 (.A1(\buffer[13][4][1] [9]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][4][1] [9]), .ZN(n_5_41_89));
   NAND4_X1 i_5_41_100 (.A1(n_5_41_98), .A2(n_5_41_96), .A3(n_5_41_94), .A4(
      n_5_41_90), .ZN(\output_filter[4][1] [10]));
   AOI221_X1 i_5_41_101 (.A(n_5_41_91), .B1(n_25), .B2(\buffer[0][4][1] [10]), 
      .C1(\buffer[12][4][1] [10]), .C2(n_27), .ZN(n_5_41_90));
   NAND4_X1 i_5_41_102 (.A1(n_5_41_97), .A2(n_5_41_95), .A3(n_5_41_93), .A4(
      n_5_41_92), .ZN(n_5_41_91));
   AOI22_X1 i_5_41_103 (.A1(\buffer[15][4][1] [10]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][1] [10]), .ZN(n_5_41_92));
   AOI22_X1 i_5_41_104 (.A1(\buffer[10][4][1] [10]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][1] [10]), .ZN(n_5_41_93));
   AOI22_X1 i_5_41_105 (.A1(\buffer[6][4][1] [10]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][4][1] [10]), .ZN(n_5_41_94));
   AOI22_X1 i_5_41_106 (.A1(\buffer[9][4][1] [10]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][4][1] [10]), .ZN(n_5_41_95));
   AOI22_X1 i_5_41_107 (.A1(\buffer[14][4][1] [10]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][1] [10]), .ZN(n_5_41_96));
   AOI22_X1 i_5_41_108 (.A1(\buffer[11][4][1] [10]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][1] [10]), .ZN(n_5_41_97));
   AOI22_X1 i_5_41_109 (.A1(\buffer[13][4][1] [10]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][1] [10]), .ZN(n_5_41_98));
   NAND4_X1 i_5_41_110 (.A1(n_5_41_107), .A2(n_5_41_105), .A3(n_5_41_103), 
      .A4(n_5_41_99), .ZN(\output_filter[4][1] [11]));
   AOI221_X1 i_5_41_111 (.A(n_5_41_100), .B1(n_25), .B2(\buffer[0][4][1] [11]), 
      .C1(\buffer[12][4][1] [11]), .C2(n_27), .ZN(n_5_41_99));
   NAND4_X1 i_5_41_112 (.A1(n_5_41_106), .A2(n_5_41_104), .A3(n_5_41_102), 
      .A4(n_5_41_101), .ZN(n_5_41_100));
   AOI22_X1 i_5_41_113 (.A1(\buffer[15][4][1] [11]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][1] [11]), .ZN(n_5_41_101));
   AOI22_X1 i_5_41_114 (.A1(\buffer[10][4][1] [11]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][1] [11]), .ZN(n_5_41_102));
   AOI22_X1 i_5_41_115 (.A1(\buffer[6][4][1] [11]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][4][1] [11]), .ZN(n_5_41_103));
   AOI22_X1 i_5_41_116 (.A1(\buffer[9][4][1] [11]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][4][1] [11]), .ZN(n_5_41_104));
   AOI22_X1 i_5_41_117 (.A1(\buffer[14][4][1] [11]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][1] [11]), .ZN(n_5_41_105));
   AOI22_X1 i_5_41_118 (.A1(\buffer[11][4][1] [11]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][1] [11]), .ZN(n_5_41_106));
   AOI22_X1 i_5_41_119 (.A1(\buffer[13][4][1] [11]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][4][1] [11]), .ZN(n_5_41_107));
   NAND4_X1 i_5_41_120 (.A1(n_5_41_116), .A2(n_5_41_114), .A3(n_5_41_112), 
      .A4(n_5_41_108), .ZN(\output_filter[4][1] [12]));
   AOI221_X1 i_5_41_121 (.A(n_5_41_109), .B1(n_25), .B2(\buffer[0][4][1] [12]), 
      .C1(\buffer[12][4][1] [12]), .C2(n_27), .ZN(n_5_41_108));
   NAND4_X1 i_5_41_122 (.A1(n_5_41_115), .A2(n_5_41_113), .A3(n_5_41_111), 
      .A4(n_5_41_110), .ZN(n_5_41_109));
   AOI22_X1 i_5_41_123 (.A1(\buffer[15][4][1] [12]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][1] [12]), .ZN(n_5_41_110));
   AOI22_X1 i_5_41_124 (.A1(\buffer[10][4][1] [12]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][1] [12]), .ZN(n_5_41_111));
   AOI22_X1 i_5_41_125 (.A1(\buffer[6][4][1] [12]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][4][1] [12]), .ZN(n_5_41_112));
   AOI22_X1 i_5_41_126 (.A1(\buffer[9][4][1] [12]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][4][1] [12]), .ZN(n_5_41_113));
   AOI22_X1 i_5_41_127 (.A1(\buffer[14][4][1] [12]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][1] [12]), .ZN(n_5_41_114));
   AOI22_X1 i_5_41_128 (.A1(\buffer[11][4][1] [12]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][1] [12]), .ZN(n_5_41_115));
   AOI22_X1 i_5_41_129 (.A1(\buffer[13][4][1] [12]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][1] [12]), .ZN(n_5_41_116));
   NAND4_X1 i_5_41_130 (.A1(n_5_41_125), .A2(n_5_41_123), .A3(n_5_41_121), 
      .A4(n_5_41_117), .ZN(\output_filter[4][1] [13]));
   AOI221_X1 i_5_41_131 (.A(n_5_41_118), .B1(n_25), .B2(\buffer[0][4][1] [13]), 
      .C1(\buffer[12][4][1] [13]), .C2(n_27), .ZN(n_5_41_117));
   NAND4_X1 i_5_41_132 (.A1(n_5_41_124), .A2(n_5_41_122), .A3(n_5_41_120), 
      .A4(n_5_41_119), .ZN(n_5_41_118));
   AOI22_X1 i_5_41_133 (.A1(\buffer[15][4][1] [13]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][1] [13]), .ZN(n_5_41_119));
   AOI22_X1 i_5_41_134 (.A1(\buffer[10][4][1] [13]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][1] [13]), .ZN(n_5_41_120));
   AOI22_X1 i_5_41_135 (.A1(\buffer[6][4][1] [13]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][4][1] [13]), .ZN(n_5_41_121));
   AOI22_X1 i_5_41_136 (.A1(\buffer[9][4][1] [13]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][4][1] [13]), .ZN(n_5_41_122));
   AOI22_X1 i_5_41_137 (.A1(\buffer[14][4][1] [13]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][1] [13]), .ZN(n_5_41_123));
   AOI22_X1 i_5_41_138 (.A1(\buffer[11][4][1] [13]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][1] [13]), .ZN(n_5_41_124));
   AOI22_X1 i_5_41_139 (.A1(\buffer[13][4][1] [13]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][4][1] [13]), .ZN(n_5_41_125));
   NAND4_X1 i_5_41_140 (.A1(n_5_41_134), .A2(n_5_41_132), .A3(n_5_41_130), 
      .A4(n_5_41_126), .ZN(\output_filter[4][1] [14]));
   AOI221_X1 i_5_41_141 (.A(n_5_41_127), .B1(n_25), .B2(\buffer[0][4][1] [14]), 
      .C1(\buffer[12][4][1] [14]), .C2(n_27), .ZN(n_5_41_126));
   NAND4_X1 i_5_41_142 (.A1(n_5_41_133), .A2(n_5_41_131), .A3(n_5_41_129), 
      .A4(n_5_41_128), .ZN(n_5_41_127));
   AOI22_X1 i_5_41_143 (.A1(\buffer[15][4][1] [14]), .A2(n_22), .B1(n_16), 
      .B2(\buffer[8][4][1] [14]), .ZN(n_5_41_128));
   AOI22_X1 i_5_41_144 (.A1(\buffer[10][4][1] [14]), .A2(n_21), .B1(n_29), 
      .B2(\buffer[7][4][1] [14]), .ZN(n_5_41_129));
   AOI22_X1 i_5_41_145 (.A1(\buffer[6][4][1] [14]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][4][1] [14]), .ZN(n_5_41_130));
   AOI22_X1 i_5_41_146 (.A1(\buffer[9][4][1] [14]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][4][1] [14]), .ZN(n_5_41_131));
   AOI22_X1 i_5_41_147 (.A1(\buffer[14][4][1] [14]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][1] [14]), .ZN(n_5_41_132));
   AOI22_X1 i_5_41_148 (.A1(\buffer[11][4][1] [14]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][1] [14]), .ZN(n_5_41_133));
   AOI22_X1 i_5_41_149 (.A1(\buffer[13][4][1] [14]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][1] [14]), .ZN(n_5_41_134));
   NAND2_X1 i_5_41_150 (.A1(n_5_41_137), .A2(n_5_41_135), .ZN(
      \output_filter[4][1] [15]));
   AOI221_X1 i_5_41_151 (.A(n_5_41_136), .B1(n_31), .B2(\buffer[3][4][1] [15]), 
      .C1(\buffer[14][4][1] [15]), .C2(n_19), .ZN(n_5_41_135));
   NAND3_X1 i_5_41_152 (.A1(n_5_41_143), .A2(n_5_41_141), .A3(n_5_41_139), 
      .ZN(n_5_41_136));
   AOI221_X1 i_5_41_153 (.A(n_5_41_138), .B1(n_16), .B2(\buffer[8][4][1] [15]), 
      .C1(\buffer[13][4][1] [15]), .C2(n_26), .ZN(n_5_41_137));
   NAND3_X1 i_5_41_154 (.A1(n_5_41_144), .A2(n_5_41_142), .A3(n_5_41_140), 
      .ZN(n_5_41_138));
   AOI22_X1 i_5_41_155 (.A1(\buffer[11][4][1] [15]), .A2(n_17), .B1(n_24), 
      .B2(\buffer[2][4][1] [15]), .ZN(n_5_41_139));
   AOI22_X1 i_5_41_156 (.A1(\buffer[10][4][1] [15]), .A2(n_21), .B1(n_23), 
      .B2(\buffer[1][4][1] [15]), .ZN(n_5_41_140));
   AOI22_X1 i_5_41_157 (.A1(\buffer[6][4][1] [15]), .A2(n_28), .B1(n_18), 
      .B2(\buffer[5][4][1] [15]), .ZN(n_5_41_141));
   AOI22_X1 i_5_41_158 (.A1(\buffer[9][4][1] [15]), .A2(n_20), .B1(n_30), 
      .B2(\buffer[4][4][1] [15]), .ZN(n_5_41_142));
   AOI22_X1 i_5_41_159 (.A1(\buffer[7][4][1] [15]), .A2(n_29), .B1(n_25), 
      .B2(\buffer[0][4][1] [15]), .ZN(n_5_41_143));
   AOI22_X1 i_5_41_160 (.A1(\buffer[15][4][1] [15]), .A2(n_22), .B1(n_27), 
      .B2(\buffer[12][4][1] [15]), .ZN(n_5_41_144));
   NAND4_X1 i_6_40_0 (.A1(n_6_40_8), .A2(n_6_40_6), .A3(n_6_40_4), .A4(n_6_40_0), 
      .ZN(\output_filter[4][0] [0]));
   AOI221_X1 i_6_40_1 (.A(n_6_40_1), .B1(n_25), .B2(\buffer[0][4][0] [0]), 
      .C1(\buffer[12][4][0] [0]), .C2(n_27), .ZN(n_6_40_0));
   NAND4_X1 i_6_40_2 (.A1(n_6_40_7), .A2(n_6_40_5), .A3(n_6_40_3), .A4(n_6_40_2), 
      .ZN(n_6_40_1));
   AOI22_X1 i_6_40_3 (.A1(\buffer[15][4][0] [0]), .A2(n_22), .B1(n_29), .B2(
      \buffer[7][4][0] [0]), .ZN(n_6_40_2));
   AOI22_X1 i_6_40_4 (.A1(\buffer[10][4][0] [0]), .A2(n_21), .B1(n_16), .B2(
      \buffer[8][4][0] [0]), .ZN(n_6_40_3));
   AOI22_X1 i_6_40_5 (.A1(\buffer[6][4][0] [0]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][0] [0]), .ZN(n_6_40_4));
   AOI22_X1 i_6_40_6 (.A1(\buffer[9][4][0] [0]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][0] [0]), .ZN(n_6_40_5));
   AOI22_X1 i_6_40_7 (.A1(\buffer[14][4][0] [0]), .A2(n_19), .B1(n_23), .B2(
      \buffer[1][4][0] [0]), .ZN(n_6_40_6));
   AOI22_X1 i_6_40_8 (.A1(\buffer[11][4][0] [0]), .A2(n_17), .B1(n_18), .B2(
      \buffer[5][4][0] [0]), .ZN(n_6_40_7));
   AOI22_X1 i_6_40_9 (.A1(\buffer[13][4][0] [0]), .A2(n_26), .B1(n_24), .B2(
      \buffer[2][4][0] [0]), .ZN(n_6_40_8));
   NAND4_X1 i_6_40_10 (.A1(n_6_40_17), .A2(n_6_40_15), .A3(n_6_40_13), .A4(
      n_6_40_9), .ZN(\output_filter[4][0] [1]));
   AOI221_X1 i_6_40_11 (.A(n_6_40_10), .B1(n_25), .B2(\buffer[0][4][0] [1]), 
      .C1(\buffer[12][4][0] [1]), .C2(n_27), .ZN(n_6_40_9));
   NAND4_X1 i_6_40_12 (.A1(n_6_40_16), .A2(n_6_40_14), .A3(n_6_40_12), .A4(
      n_6_40_11), .ZN(n_6_40_10));
   AOI22_X1 i_6_40_13 (.A1(\buffer[15][4][0] [1]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][0] [1]), .ZN(n_6_40_11));
   AOI22_X1 i_6_40_14 (.A1(\buffer[10][4][0] [1]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][0] [1]), .ZN(n_6_40_12));
   AOI22_X1 i_6_40_15 (.A1(\buffer[6][4][0] [1]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][0] [1]), .ZN(n_6_40_13));
   AOI22_X1 i_6_40_16 (.A1(\buffer[9][4][0] [1]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][0] [1]), .ZN(n_6_40_14));
   AOI22_X1 i_6_40_17 (.A1(\buffer[14][4][0] [1]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][0] [1]), .ZN(n_6_40_15));
   AOI22_X1 i_6_40_18 (.A1(\buffer[11][4][0] [1]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][0] [1]), .ZN(n_6_40_16));
   AOI22_X1 i_6_40_19 (.A1(\buffer[13][4][0] [1]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][0] [1]), .ZN(n_6_40_17));
   NAND4_X1 i_6_40_20 (.A1(n_6_40_26), .A2(n_6_40_24), .A3(n_6_40_22), .A4(
      n_6_40_18), .ZN(\output_filter[4][0] [2]));
   AOI221_X1 i_6_40_21 (.A(n_6_40_19), .B1(n_25), .B2(\buffer[0][4][0] [2]), 
      .C1(\buffer[12][4][0] [2]), .C2(n_27), .ZN(n_6_40_18));
   NAND4_X1 i_6_40_22 (.A1(n_6_40_25), .A2(n_6_40_23), .A3(n_6_40_21), .A4(
      n_6_40_20), .ZN(n_6_40_19));
   AOI22_X1 i_6_40_23 (.A1(\buffer[15][4][0] [2]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][0] [2]), .ZN(n_6_40_20));
   AOI22_X1 i_6_40_24 (.A1(\buffer[10][4][0] [2]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][0] [2]), .ZN(n_6_40_21));
   AOI22_X1 i_6_40_25 (.A1(\buffer[6][4][0] [2]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][0] [2]), .ZN(n_6_40_22));
   AOI22_X1 i_6_40_26 (.A1(\buffer[9][4][0] [2]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][0] [2]), .ZN(n_6_40_23));
   AOI22_X1 i_6_40_27 (.A1(\buffer[14][4][0] [2]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][0] [2]), .ZN(n_6_40_24));
   AOI22_X1 i_6_40_28 (.A1(\buffer[11][4][0] [2]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][0] [2]), .ZN(n_6_40_25));
   AOI22_X1 i_6_40_29 (.A1(\buffer[13][4][0] [2]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][0] [2]), .ZN(n_6_40_26));
   NAND4_X1 i_6_40_30 (.A1(n_6_40_35), .A2(n_6_40_33), .A3(n_6_40_31), .A4(
      n_6_40_27), .ZN(\output_filter[4][0] [3]));
   AOI221_X1 i_6_40_31 (.A(n_6_40_28), .B1(n_25), .B2(\buffer[0][4][0] [3]), 
      .C1(\buffer[12][4][0] [3]), .C2(n_27), .ZN(n_6_40_27));
   NAND4_X1 i_6_40_32 (.A1(n_6_40_34), .A2(n_6_40_32), .A3(n_6_40_30), .A4(
      n_6_40_29), .ZN(n_6_40_28));
   AOI22_X1 i_6_40_33 (.A1(\buffer[15][4][0] [3]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][0] [3]), .ZN(n_6_40_29));
   AOI22_X1 i_6_40_34 (.A1(\buffer[10][4][0] [3]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][0] [3]), .ZN(n_6_40_30));
   AOI22_X1 i_6_40_35 (.A1(\buffer[6][4][0] [3]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][0] [3]), .ZN(n_6_40_31));
   AOI22_X1 i_6_40_36 (.A1(\buffer[9][4][0] [3]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][0] [3]), .ZN(n_6_40_32));
   AOI22_X1 i_6_40_37 (.A1(\buffer[14][4][0] [3]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][0] [3]), .ZN(n_6_40_33));
   AOI22_X1 i_6_40_38 (.A1(\buffer[11][4][0] [3]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][0] [3]), .ZN(n_6_40_34));
   AOI22_X1 i_6_40_39 (.A1(\buffer[13][4][0] [3]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][0] [3]), .ZN(n_6_40_35));
   NAND4_X1 i_6_40_40 (.A1(n_6_40_44), .A2(n_6_40_42), .A3(n_6_40_40), .A4(
      n_6_40_36), .ZN(\output_filter[4][0] [4]));
   AOI221_X1 i_6_40_41 (.A(n_6_40_37), .B1(n_25), .B2(\buffer[0][4][0] [4]), 
      .C1(\buffer[12][4][0] [4]), .C2(n_27), .ZN(n_6_40_36));
   NAND4_X1 i_6_40_42 (.A1(n_6_40_43), .A2(n_6_40_41), .A3(n_6_40_39), .A4(
      n_6_40_38), .ZN(n_6_40_37));
   AOI22_X1 i_6_40_43 (.A1(\buffer[15][4][0] [4]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][0] [4]), .ZN(n_6_40_38));
   AOI22_X1 i_6_40_44 (.A1(\buffer[10][4][0] [4]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][0] [4]), .ZN(n_6_40_39));
   AOI22_X1 i_6_40_45 (.A1(\buffer[6][4][0] [4]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][0] [4]), .ZN(n_6_40_40));
   AOI22_X1 i_6_40_46 (.A1(\buffer[9][4][0] [4]), .A2(n_20), .B1(n_24), .B2(
      \buffer[2][4][0] [4]), .ZN(n_6_40_41));
   AOI22_X1 i_6_40_47 (.A1(\buffer[14][4][0] [4]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][0] [4]), .ZN(n_6_40_42));
   AOI22_X1 i_6_40_48 (.A1(\buffer[11][4][0] [4]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][0] [4]), .ZN(n_6_40_43));
   AOI22_X1 i_6_40_49 (.A1(\buffer[13][4][0] [4]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][4][0] [4]), .ZN(n_6_40_44));
   NAND4_X1 i_6_40_50 (.A1(n_6_40_53), .A2(n_6_40_51), .A3(n_6_40_49), .A4(
      n_6_40_45), .ZN(\output_filter[4][0] [5]));
   AOI221_X1 i_6_40_51 (.A(n_6_40_46), .B1(n_25), .B2(\buffer[0][4][0] [5]), 
      .C1(\buffer[12][4][0] [5]), .C2(n_27), .ZN(n_6_40_45));
   NAND4_X1 i_6_40_52 (.A1(n_6_40_52), .A2(n_6_40_50), .A3(n_6_40_48), .A4(
      n_6_40_47), .ZN(n_6_40_46));
   AOI22_X1 i_6_40_53 (.A1(\buffer[15][4][0] [5]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][0] [5]), .ZN(n_6_40_47));
   AOI22_X1 i_6_40_54 (.A1(\buffer[10][4][0] [5]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][0] [5]), .ZN(n_6_40_48));
   AOI22_X1 i_6_40_55 (.A1(\buffer[6][4][0] [5]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][0] [5]), .ZN(n_6_40_49));
   AOI22_X1 i_6_40_56 (.A1(\buffer[9][4][0] [5]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][0] [5]), .ZN(n_6_40_50));
   AOI22_X1 i_6_40_57 (.A1(\buffer[14][4][0] [5]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][0] [5]), .ZN(n_6_40_51));
   AOI22_X1 i_6_40_58 (.A1(\buffer[11][4][0] [5]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][0] [5]), .ZN(n_6_40_52));
   AOI22_X1 i_6_40_59 (.A1(\buffer[13][4][0] [5]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][0] [5]), .ZN(n_6_40_53));
   NAND4_X1 i_6_40_60 (.A1(n_6_40_62), .A2(n_6_40_60), .A3(n_6_40_58), .A4(
      n_6_40_54), .ZN(\output_filter[4][0] [6]));
   AOI221_X1 i_6_40_61 (.A(n_6_40_55), .B1(n_25), .B2(\buffer[0][4][0] [6]), 
      .C1(\buffer[12][4][0] [6]), .C2(n_27), .ZN(n_6_40_54));
   NAND4_X1 i_6_40_62 (.A1(n_6_40_61), .A2(n_6_40_59), .A3(n_6_40_57), .A4(
      n_6_40_56), .ZN(n_6_40_55));
   AOI22_X1 i_6_40_63 (.A1(\buffer[15][4][0] [6]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][0] [6]), .ZN(n_6_40_56));
   AOI22_X1 i_6_40_64 (.A1(\buffer[10][4][0] [6]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][0] [6]), .ZN(n_6_40_57));
   AOI22_X1 i_6_40_65 (.A1(\buffer[6][4][0] [6]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][0] [6]), .ZN(n_6_40_58));
   AOI22_X1 i_6_40_66 (.A1(\buffer[9][4][0] [6]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][0] [6]), .ZN(n_6_40_59));
   AOI22_X1 i_6_40_67 (.A1(\buffer[14][4][0] [6]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][0] [6]), .ZN(n_6_40_60));
   AOI22_X1 i_6_40_68 (.A1(\buffer[11][4][0] [6]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][0] [6]), .ZN(n_6_40_61));
   AOI22_X1 i_6_40_69 (.A1(\buffer[13][4][0] [6]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][0] [6]), .ZN(n_6_40_62));
   NAND4_X1 i_6_40_70 (.A1(n_6_40_71), .A2(n_6_40_69), .A3(n_6_40_67), .A4(
      n_6_40_63), .ZN(\output_filter[4][0] [7]));
   AOI221_X1 i_6_40_71 (.A(n_6_40_64), .B1(n_25), .B2(\buffer[0][4][0] [7]), 
      .C1(\buffer[12][4][0] [7]), .C2(n_27), .ZN(n_6_40_63));
   NAND4_X1 i_6_40_72 (.A1(n_6_40_70), .A2(n_6_40_68), .A3(n_6_40_66), .A4(
      n_6_40_65), .ZN(n_6_40_64));
   AOI22_X1 i_6_40_73 (.A1(\buffer[15][4][0] [7]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][0] [7]), .ZN(n_6_40_65));
   AOI22_X1 i_6_40_74 (.A1(\buffer[10][4][0] [7]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][0] [7]), .ZN(n_6_40_66));
   AOI22_X1 i_6_40_75 (.A1(\buffer[6][4][0] [7]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][0] [7]), .ZN(n_6_40_67));
   AOI22_X1 i_6_40_76 (.A1(\buffer[9][4][0] [7]), .A2(n_20), .B1(n_24), .B2(
      \buffer[2][4][0] [7]), .ZN(n_6_40_68));
   AOI22_X1 i_6_40_77 (.A1(\buffer[14][4][0] [7]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][0] [7]), .ZN(n_6_40_69));
   AOI22_X1 i_6_40_78 (.A1(\buffer[11][4][0] [7]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][0] [7]), .ZN(n_6_40_70));
   AOI22_X1 i_6_40_79 (.A1(\buffer[13][4][0] [7]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][4][0] [7]), .ZN(n_6_40_71));
   NAND4_X1 i_6_40_80 (.A1(n_6_40_80), .A2(n_6_40_78), .A3(n_6_40_76), .A4(
      n_6_40_72), .ZN(\output_filter[4][0] [8]));
   AOI221_X1 i_6_40_81 (.A(n_6_40_73), .B1(n_25), .B2(\buffer[0][4][0] [8]), 
      .C1(\buffer[12][4][0] [8]), .C2(n_27), .ZN(n_6_40_72));
   NAND4_X1 i_6_40_82 (.A1(n_6_40_79), .A2(n_6_40_77), .A3(n_6_40_75), .A4(
      n_6_40_74), .ZN(n_6_40_73));
   AOI22_X1 i_6_40_83 (.A1(\buffer[15][4][0] [8]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][0] [8]), .ZN(n_6_40_74));
   AOI22_X1 i_6_40_84 (.A1(\buffer[10][4][0] [8]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][0] [8]), .ZN(n_6_40_75));
   AOI22_X1 i_6_40_85 (.A1(\buffer[6][4][0] [8]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][0] [8]), .ZN(n_6_40_76));
   AOI22_X1 i_6_40_86 (.A1(\buffer[9][4][0] [8]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][4][0] [8]), .ZN(n_6_40_77));
   AOI22_X1 i_6_40_87 (.A1(\buffer[14][4][0] [8]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][0] [8]), .ZN(n_6_40_78));
   AOI22_X1 i_6_40_88 (.A1(\buffer[11][4][0] [8]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][0] [8]), .ZN(n_6_40_79));
   AOI22_X1 i_6_40_89 (.A1(\buffer[13][4][0] [8]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][0] [8]), .ZN(n_6_40_80));
   NAND4_X1 i_6_40_90 (.A1(n_6_40_89), .A2(n_6_40_87), .A3(n_6_40_85), .A4(
      n_6_40_81), .ZN(\output_filter[4][0] [9]));
   AOI221_X1 i_6_40_91 (.A(n_6_40_82), .B1(n_25), .B2(\buffer[0][4][0] [9]), 
      .C1(\buffer[12][4][0] [9]), .C2(n_27), .ZN(n_6_40_81));
   NAND4_X1 i_6_40_92 (.A1(n_6_40_88), .A2(n_6_40_86), .A3(n_6_40_84), .A4(
      n_6_40_83), .ZN(n_6_40_82));
   AOI22_X1 i_6_40_93 (.A1(\buffer[15][4][0] [9]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][0] [9]), .ZN(n_6_40_83));
   AOI22_X1 i_6_40_94 (.A1(\buffer[10][4][0] [9]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][0] [9]), .ZN(n_6_40_84));
   AOI22_X1 i_6_40_95 (.A1(\buffer[6][4][0] [9]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][4][0] [9]), .ZN(n_6_40_85));
   AOI22_X1 i_6_40_96 (.A1(\buffer[9][4][0] [9]), .A2(n_20), .B1(n_24), .B2(
      \buffer[2][4][0] [9]), .ZN(n_6_40_86));
   AOI22_X1 i_6_40_97 (.A1(\buffer[14][4][0] [9]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][0] [9]), .ZN(n_6_40_87));
   AOI22_X1 i_6_40_98 (.A1(\buffer[11][4][0] [9]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][0] [9]), .ZN(n_6_40_88));
   AOI22_X1 i_6_40_99 (.A1(\buffer[13][4][0] [9]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][4][0] [9]), .ZN(n_6_40_89));
   NAND4_X1 i_6_40_100 (.A1(n_6_40_98), .A2(n_6_40_96), .A3(n_6_40_94), .A4(
      n_6_40_90), .ZN(\output_filter[4][0] [10]));
   AOI221_X1 i_6_40_101 (.A(n_6_40_91), .B1(n_25), .B2(\buffer[0][4][0] [10]), 
      .C1(\buffer[12][4][0] [10]), .C2(n_27), .ZN(n_6_40_90));
   NAND4_X1 i_6_40_102 (.A1(n_6_40_97), .A2(n_6_40_95), .A3(n_6_40_93), .A4(
      n_6_40_92), .ZN(n_6_40_91));
   AOI22_X1 i_6_40_103 (.A1(\buffer[15][4][0] [10]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][0] [10]), .ZN(n_6_40_92));
   AOI22_X1 i_6_40_104 (.A1(\buffer[10][4][0] [10]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][0] [10]), .ZN(n_6_40_93));
   AOI22_X1 i_6_40_105 (.A1(\buffer[6][4][0] [10]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][4][0] [10]), .ZN(n_6_40_94));
   AOI22_X1 i_6_40_106 (.A1(\buffer[9][4][0] [10]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][4][0] [10]), .ZN(n_6_40_95));
   AOI22_X1 i_6_40_107 (.A1(\buffer[14][4][0] [10]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][0] [10]), .ZN(n_6_40_96));
   AOI22_X1 i_6_40_108 (.A1(\buffer[11][4][0] [10]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][0] [10]), .ZN(n_6_40_97));
   AOI22_X1 i_6_40_109 (.A1(\buffer[13][4][0] [10]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][0] [10]), .ZN(n_6_40_98));
   NAND4_X1 i_6_40_110 (.A1(n_6_40_107), .A2(n_6_40_105), .A3(n_6_40_103), 
      .A4(n_6_40_99), .ZN(\output_filter[4][0] [11]));
   AOI221_X1 i_6_40_111 (.A(n_6_40_100), .B1(n_25), .B2(\buffer[0][4][0] [11]), 
      .C1(\buffer[12][4][0] [11]), .C2(n_27), .ZN(n_6_40_99));
   NAND4_X1 i_6_40_112 (.A1(n_6_40_106), .A2(n_6_40_104), .A3(n_6_40_102), 
      .A4(n_6_40_101), .ZN(n_6_40_100));
   AOI22_X1 i_6_40_113 (.A1(\buffer[15][4][0] [11]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][0] [11]), .ZN(n_6_40_101));
   AOI22_X1 i_6_40_114 (.A1(\buffer[10][4][0] [11]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][0] [11]), .ZN(n_6_40_102));
   AOI22_X1 i_6_40_115 (.A1(\buffer[6][4][0] [11]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][4][0] [11]), .ZN(n_6_40_103));
   AOI22_X1 i_6_40_116 (.A1(\buffer[9][4][0] [11]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][4][0] [11]), .ZN(n_6_40_104));
   AOI22_X1 i_6_40_117 (.A1(\buffer[14][4][0] [11]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][0] [11]), .ZN(n_6_40_105));
   AOI22_X1 i_6_40_118 (.A1(\buffer[11][4][0] [11]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][0] [11]), .ZN(n_6_40_106));
   AOI22_X1 i_6_40_119 (.A1(\buffer[13][4][0] [11]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][4][0] [11]), .ZN(n_6_40_107));
   NAND4_X1 i_6_40_120 (.A1(n_6_40_116), .A2(n_6_40_114), .A3(n_6_40_112), 
      .A4(n_6_40_108), .ZN(\output_filter[4][0] [12]));
   AOI221_X1 i_6_40_121 (.A(n_6_40_109), .B1(n_25), .B2(\buffer[0][4][0] [12]), 
      .C1(\buffer[12][4][0] [12]), .C2(n_27), .ZN(n_6_40_108));
   NAND4_X1 i_6_40_122 (.A1(n_6_40_115), .A2(n_6_40_113), .A3(n_6_40_111), 
      .A4(n_6_40_110), .ZN(n_6_40_109));
   AOI22_X1 i_6_40_123 (.A1(\buffer[15][4][0] [12]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][0] [12]), .ZN(n_6_40_110));
   AOI22_X1 i_6_40_124 (.A1(\buffer[10][4][0] [12]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][0] [12]), .ZN(n_6_40_111));
   AOI22_X1 i_6_40_125 (.A1(\buffer[6][4][0] [12]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][4][0] [12]), .ZN(n_6_40_112));
   AOI22_X1 i_6_40_126 (.A1(\buffer[9][4][0] [12]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][4][0] [12]), .ZN(n_6_40_113));
   AOI22_X1 i_6_40_127 (.A1(\buffer[14][4][0] [12]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][0] [12]), .ZN(n_6_40_114));
   AOI22_X1 i_6_40_128 (.A1(\buffer[11][4][0] [12]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][0] [12]), .ZN(n_6_40_115));
   AOI22_X1 i_6_40_129 (.A1(\buffer[13][4][0] [12]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][0] [12]), .ZN(n_6_40_116));
   NAND4_X1 i_6_40_130 (.A1(n_6_40_125), .A2(n_6_40_123), .A3(n_6_40_121), 
      .A4(n_6_40_117), .ZN(\output_filter[4][0] [13]));
   AOI221_X1 i_6_40_131 (.A(n_6_40_118), .B1(n_25), .B2(\buffer[0][4][0] [13]), 
      .C1(\buffer[12][4][0] [13]), .C2(n_27), .ZN(n_6_40_117));
   NAND4_X1 i_6_40_132 (.A1(n_6_40_124), .A2(n_6_40_122), .A3(n_6_40_120), 
      .A4(n_6_40_119), .ZN(n_6_40_118));
   AOI22_X1 i_6_40_133 (.A1(\buffer[15][4][0] [13]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][4][0] [13]), .ZN(n_6_40_119));
   AOI22_X1 i_6_40_134 (.A1(\buffer[10][4][0] [13]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][4][0] [13]), .ZN(n_6_40_120));
   AOI22_X1 i_6_40_135 (.A1(\buffer[6][4][0] [13]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][4][0] [13]), .ZN(n_6_40_121));
   AOI22_X1 i_6_40_136 (.A1(\buffer[9][4][0] [13]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][4][0] [13]), .ZN(n_6_40_122));
   AOI22_X1 i_6_40_137 (.A1(\buffer[14][4][0] [13]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][0] [13]), .ZN(n_6_40_123));
   AOI22_X1 i_6_40_138 (.A1(\buffer[11][4][0] [13]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][0] [13]), .ZN(n_6_40_124));
   AOI22_X1 i_6_40_139 (.A1(\buffer[13][4][0] [13]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][4][0] [13]), .ZN(n_6_40_125));
   NAND4_X1 i_6_40_140 (.A1(n_6_40_134), .A2(n_6_40_132), .A3(n_6_40_130), 
      .A4(n_6_40_126), .ZN(\output_filter[4][0] [14]));
   AOI221_X1 i_6_40_141 (.A(n_6_40_127), .B1(n_25), .B2(\buffer[0][4][0] [14]), 
      .C1(\buffer[12][4][0] [14]), .C2(n_27), .ZN(n_6_40_126));
   NAND4_X1 i_6_40_142 (.A1(n_6_40_133), .A2(n_6_40_131), .A3(n_6_40_129), 
      .A4(n_6_40_128), .ZN(n_6_40_127));
   AOI22_X1 i_6_40_143 (.A1(\buffer[15][4][0] [14]), .A2(n_22), .B1(n_16), 
      .B2(\buffer[8][4][0] [14]), .ZN(n_6_40_128));
   AOI22_X1 i_6_40_144 (.A1(\buffer[10][4][0] [14]), .A2(n_21), .B1(n_29), 
      .B2(\buffer[7][4][0] [14]), .ZN(n_6_40_129));
   AOI22_X1 i_6_40_145 (.A1(\buffer[6][4][0] [14]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][4][0] [14]), .ZN(n_6_40_130));
   AOI22_X1 i_6_40_146 (.A1(\buffer[9][4][0] [14]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][4][0] [14]), .ZN(n_6_40_131));
   AOI22_X1 i_6_40_147 (.A1(\buffer[14][4][0] [14]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][4][0] [14]), .ZN(n_6_40_132));
   AOI22_X1 i_6_40_148 (.A1(\buffer[11][4][0] [14]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][4][0] [14]), .ZN(n_6_40_133));
   AOI22_X1 i_6_40_149 (.A1(\buffer[13][4][0] [14]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][4][0] [14]), .ZN(n_6_40_134));
   NAND2_X1 i_6_40_150 (.A1(n_6_40_137), .A2(n_6_40_135), .ZN(
      \output_filter[4][0] [15]));
   AOI221_X1 i_6_40_151 (.A(n_6_40_136), .B1(n_31), .B2(\buffer[3][4][0] [15]), 
      .C1(\buffer[14][4][0] [15]), .C2(n_19), .ZN(n_6_40_135));
   NAND3_X1 i_6_40_152 (.A1(n_6_40_143), .A2(n_6_40_141), .A3(n_6_40_139), 
      .ZN(n_6_40_136));
   AOI221_X1 i_6_40_153 (.A(n_6_40_138), .B1(n_16), .B2(\buffer[8][4][0] [15]), 
      .C1(\buffer[13][4][0] [15]), .C2(n_26), .ZN(n_6_40_137));
   NAND3_X1 i_6_40_154 (.A1(n_6_40_144), .A2(n_6_40_142), .A3(n_6_40_140), 
      .ZN(n_6_40_138));
   AOI22_X1 i_6_40_155 (.A1(\buffer[11][4][0] [15]), .A2(n_17), .B1(n_24), 
      .B2(\buffer[2][4][0] [15]), .ZN(n_6_40_139));
   AOI22_X1 i_6_40_156 (.A1(\buffer[10][4][0] [15]), .A2(n_21), .B1(n_23), 
      .B2(\buffer[1][4][0] [15]), .ZN(n_6_40_140));
   AOI22_X1 i_6_40_157 (.A1(\buffer[6][4][0] [15]), .A2(n_28), .B1(n_18), 
      .B2(\buffer[5][4][0] [15]), .ZN(n_6_40_141));
   AOI22_X1 i_6_40_158 (.A1(\buffer[9][4][0] [15]), .A2(n_20), .B1(n_30), 
      .B2(\buffer[4][4][0] [15]), .ZN(n_6_40_142));
   AOI22_X1 i_6_40_159 (.A1(\buffer[7][4][0] [15]), .A2(n_29), .B1(n_25), 
      .B2(\buffer[0][4][0] [15]), .ZN(n_6_40_143));
   AOI22_X1 i_6_40_160 (.A1(\buffer[15][4][0] [15]), .A2(n_22), .B1(n_27), 
      .B2(\buffer[12][4][0] [15]), .ZN(n_6_40_144));
   NAND4_X1 i_7_39_0 (.A1(n_7_39_8), .A2(n_7_39_6), .A3(n_7_39_4), .A4(n_7_39_0), 
      .ZN(\output_filter[3][4] [0]));
   AOI221_X1 i_7_39_1 (.A(n_7_39_1), .B1(n_25), .B2(\buffer[0][3][4] [0]), 
      .C1(\buffer[12][3][4] [0]), .C2(n_27), .ZN(n_7_39_0));
   NAND4_X1 i_7_39_2 (.A1(n_7_39_7), .A2(n_7_39_5), .A3(n_7_39_3), .A4(n_7_39_2), 
      .ZN(n_7_39_1));
   AOI22_X1 i_7_39_3 (.A1(\buffer[15][3][4] [0]), .A2(n_22), .B1(n_29), .B2(
      \buffer[7][3][4] [0]), .ZN(n_7_39_2));
   AOI22_X1 i_7_39_4 (.A1(\buffer[10][3][4] [0]), .A2(n_21), .B1(n_16), .B2(
      \buffer[8][3][4] [0]), .ZN(n_7_39_3));
   AOI22_X1 i_7_39_5 (.A1(\buffer[6][3][4] [0]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][4] [0]), .ZN(n_7_39_4));
   AOI22_X1 i_7_39_6 (.A1(\buffer[9][3][4] [0]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][3][4] [0]), .ZN(n_7_39_5));
   AOI22_X1 i_7_39_7 (.A1(\buffer[14][3][4] [0]), .A2(n_19), .B1(n_23), .B2(
      \buffer[1][3][4] [0]), .ZN(n_7_39_6));
   AOI22_X1 i_7_39_8 (.A1(\buffer[11][3][4] [0]), .A2(n_17), .B1(n_18), .B2(
      \buffer[5][3][4] [0]), .ZN(n_7_39_7));
   AOI22_X1 i_7_39_9 (.A1(\buffer[13][3][4] [0]), .A2(n_26), .B1(n_24), .B2(
      \buffer[2][3][4] [0]), .ZN(n_7_39_8));
   NAND4_X1 i_7_39_10 (.A1(n_7_39_17), .A2(n_7_39_15), .A3(n_7_39_13), .A4(
      n_7_39_9), .ZN(\output_filter[3][4] [1]));
   AOI221_X1 i_7_39_11 (.A(n_7_39_10), .B1(n_25), .B2(\buffer[0][3][4] [1]), 
      .C1(\buffer[12][3][4] [1]), .C2(n_27), .ZN(n_7_39_9));
   NAND4_X1 i_7_39_12 (.A1(n_7_39_16), .A2(n_7_39_14), .A3(n_7_39_12), .A4(
      n_7_39_11), .ZN(n_7_39_10));
   AOI22_X1 i_7_39_13 (.A1(\buffer[15][3][4] [1]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][4] [1]), .ZN(n_7_39_11));
   AOI22_X1 i_7_39_14 (.A1(\buffer[10][3][4] [1]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][4] [1]), .ZN(n_7_39_12));
   AOI22_X1 i_7_39_15 (.A1(\buffer[6][3][4] [1]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][4] [1]), .ZN(n_7_39_13));
   AOI22_X1 i_7_39_16 (.A1(\buffer[9][3][4] [1]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][3][4] [1]), .ZN(n_7_39_14));
   AOI22_X1 i_7_39_17 (.A1(\buffer[14][3][4] [1]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][4] [1]), .ZN(n_7_39_15));
   AOI22_X1 i_7_39_18 (.A1(\buffer[11][3][4] [1]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][4] [1]), .ZN(n_7_39_16));
   AOI22_X1 i_7_39_19 (.A1(\buffer[13][3][4] [1]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][4] [1]), .ZN(n_7_39_17));
   NAND4_X1 i_7_39_20 (.A1(n_7_39_26), .A2(n_7_39_24), .A3(n_7_39_22), .A4(
      n_7_39_18), .ZN(\output_filter[3][4] [2]));
   AOI221_X1 i_7_39_21 (.A(n_7_39_19), .B1(n_25), .B2(\buffer[0][3][4] [2]), 
      .C1(\buffer[12][3][4] [2]), .C2(n_27), .ZN(n_7_39_18));
   NAND4_X1 i_7_39_22 (.A1(n_7_39_25), .A2(n_7_39_23), .A3(n_7_39_21), .A4(
      n_7_39_20), .ZN(n_7_39_19));
   AOI22_X1 i_7_39_23 (.A1(\buffer[15][3][4] [2]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][4] [2]), .ZN(n_7_39_20));
   AOI22_X1 i_7_39_24 (.A1(\buffer[10][3][4] [2]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][4] [2]), .ZN(n_7_39_21));
   AOI22_X1 i_7_39_25 (.A1(\buffer[6][3][4] [2]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][4] [2]), .ZN(n_7_39_22));
   AOI22_X1 i_7_39_26 (.A1(\buffer[9][3][4] [2]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][3][4] [2]), .ZN(n_7_39_23));
   AOI22_X1 i_7_39_27 (.A1(\buffer[14][3][4] [2]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][4] [2]), .ZN(n_7_39_24));
   AOI22_X1 i_7_39_28 (.A1(\buffer[11][3][4] [2]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][4] [2]), .ZN(n_7_39_25));
   AOI22_X1 i_7_39_29 (.A1(\buffer[13][3][4] [2]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][4] [2]), .ZN(n_7_39_26));
   NAND4_X1 i_7_39_30 (.A1(n_7_39_35), .A2(n_7_39_33), .A3(n_7_39_31), .A4(
      n_7_39_27), .ZN(\output_filter[3][4] [3]));
   AOI221_X1 i_7_39_31 (.A(n_7_39_28), .B1(n_25), .B2(\buffer[0][3][4] [3]), 
      .C1(\buffer[12][3][4] [3]), .C2(n_27), .ZN(n_7_39_27));
   NAND4_X1 i_7_39_32 (.A1(n_7_39_34), .A2(n_7_39_32), .A3(n_7_39_30), .A4(
      n_7_39_29), .ZN(n_7_39_28));
   AOI22_X1 i_7_39_33 (.A1(\buffer[15][3][4] [3]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][4] [3]), .ZN(n_7_39_29));
   AOI22_X1 i_7_39_34 (.A1(\buffer[10][3][4] [3]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][4] [3]), .ZN(n_7_39_30));
   AOI22_X1 i_7_39_35 (.A1(\buffer[6][3][4] [3]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][4] [3]), .ZN(n_7_39_31));
   AOI22_X1 i_7_39_36 (.A1(\buffer[9][3][4] [3]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][3][4] [3]), .ZN(n_7_39_32));
   AOI22_X1 i_7_39_37 (.A1(\buffer[14][3][4] [3]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][4] [3]), .ZN(n_7_39_33));
   AOI22_X1 i_7_39_38 (.A1(\buffer[11][3][4] [3]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][4] [3]), .ZN(n_7_39_34));
   AOI22_X1 i_7_39_39 (.A1(\buffer[13][3][4] [3]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][4] [3]), .ZN(n_7_39_35));
   NAND4_X1 i_7_39_40 (.A1(n_7_39_44), .A2(n_7_39_42), .A3(n_7_39_40), .A4(
      n_7_39_36), .ZN(\output_filter[3][4] [4]));
   AOI221_X1 i_7_39_41 (.A(n_7_39_37), .B1(n_25), .B2(\buffer[0][3][4] [4]), 
      .C1(\buffer[12][3][4] [4]), .C2(n_27), .ZN(n_7_39_36));
   NAND4_X1 i_7_39_42 (.A1(n_7_39_43), .A2(n_7_39_41), .A3(n_7_39_39), .A4(
      n_7_39_38), .ZN(n_7_39_37));
   AOI22_X1 i_7_39_43 (.A1(\buffer[15][3][4] [4]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][4] [4]), .ZN(n_7_39_38));
   AOI22_X1 i_7_39_44 (.A1(\buffer[10][3][4] [4]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][4] [4]), .ZN(n_7_39_39));
   AOI22_X1 i_7_39_45 (.A1(\buffer[6][3][4] [4]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][4] [4]), .ZN(n_7_39_40));
   AOI22_X1 i_7_39_46 (.A1(\buffer[9][3][4] [4]), .A2(n_20), .B1(n_24), .B2(
      \buffer[2][3][4] [4]), .ZN(n_7_39_41));
   AOI22_X1 i_7_39_47 (.A1(\buffer[14][3][4] [4]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][4] [4]), .ZN(n_7_39_42));
   AOI22_X1 i_7_39_48 (.A1(\buffer[11][3][4] [4]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][4] [4]), .ZN(n_7_39_43));
   AOI22_X1 i_7_39_49 (.A1(\buffer[13][3][4] [4]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][3][4] [4]), .ZN(n_7_39_44));
   NAND4_X1 i_7_39_50 (.A1(n_7_39_53), .A2(n_7_39_51), .A3(n_7_39_49), .A4(
      n_7_39_45), .ZN(\output_filter[3][4] [5]));
   AOI221_X1 i_7_39_51 (.A(n_7_39_46), .B1(n_25), .B2(\buffer[0][3][4] [5]), 
      .C1(\buffer[12][3][4] [5]), .C2(n_27), .ZN(n_7_39_45));
   NAND4_X1 i_7_39_52 (.A1(n_7_39_52), .A2(n_7_39_50), .A3(n_7_39_48), .A4(
      n_7_39_47), .ZN(n_7_39_46));
   AOI22_X1 i_7_39_53 (.A1(\buffer[15][3][4] [5]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][4] [5]), .ZN(n_7_39_47));
   AOI22_X1 i_7_39_54 (.A1(\buffer[10][3][4] [5]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][4] [5]), .ZN(n_7_39_48));
   AOI22_X1 i_7_39_55 (.A1(\buffer[6][3][4] [5]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][4] [5]), .ZN(n_7_39_49));
   AOI22_X1 i_7_39_56 (.A1(\buffer[9][3][4] [5]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][3][4] [5]), .ZN(n_7_39_50));
   AOI22_X1 i_7_39_57 (.A1(\buffer[14][3][4] [5]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][4] [5]), .ZN(n_7_39_51));
   AOI22_X1 i_7_39_58 (.A1(\buffer[11][3][4] [5]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][4] [5]), .ZN(n_7_39_52));
   AOI22_X1 i_7_39_59 (.A1(\buffer[13][3][4] [5]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][4] [5]), .ZN(n_7_39_53));
   NAND4_X1 i_7_39_60 (.A1(n_7_39_62), .A2(n_7_39_60), .A3(n_7_39_58), .A4(
      n_7_39_54), .ZN(\output_filter[3][4] [6]));
   AOI221_X1 i_7_39_61 (.A(n_7_39_55), .B1(n_25), .B2(\buffer[0][3][4] [6]), 
      .C1(\buffer[12][3][4] [6]), .C2(n_27), .ZN(n_7_39_54));
   NAND4_X1 i_7_39_62 (.A1(n_7_39_61), .A2(n_7_39_59), .A3(n_7_39_57), .A4(
      n_7_39_56), .ZN(n_7_39_55));
   AOI22_X1 i_7_39_63 (.A1(\buffer[15][3][4] [6]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][4] [6]), .ZN(n_7_39_56));
   AOI22_X1 i_7_39_64 (.A1(\buffer[10][3][4] [6]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][4] [6]), .ZN(n_7_39_57));
   AOI22_X1 i_7_39_65 (.A1(\buffer[6][3][4] [6]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][4] [6]), .ZN(n_7_39_58));
   AOI22_X1 i_7_39_66 (.A1(\buffer[9][3][4] [6]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][3][4] [6]), .ZN(n_7_39_59));
   AOI22_X1 i_7_39_67 (.A1(\buffer[14][3][4] [6]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][4] [6]), .ZN(n_7_39_60));
   AOI22_X1 i_7_39_68 (.A1(\buffer[11][3][4] [6]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][4] [6]), .ZN(n_7_39_61));
   AOI22_X1 i_7_39_69 (.A1(\buffer[13][3][4] [6]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][4] [6]), .ZN(n_7_39_62));
   NAND4_X1 i_7_39_70 (.A1(n_7_39_71), .A2(n_7_39_69), .A3(n_7_39_67), .A4(
      n_7_39_63), .ZN(\output_filter[3][4] [7]));
   AOI221_X1 i_7_39_71 (.A(n_7_39_64), .B1(n_25), .B2(\buffer[0][3][4] [7]), 
      .C1(\buffer[12][3][4] [7]), .C2(n_27), .ZN(n_7_39_63));
   NAND4_X1 i_7_39_72 (.A1(n_7_39_70), .A2(n_7_39_68), .A3(n_7_39_66), .A4(
      n_7_39_65), .ZN(n_7_39_64));
   AOI22_X1 i_7_39_73 (.A1(\buffer[15][3][4] [7]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][4] [7]), .ZN(n_7_39_65));
   AOI22_X1 i_7_39_74 (.A1(\buffer[10][3][4] [7]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][4] [7]), .ZN(n_7_39_66));
   AOI22_X1 i_7_39_75 (.A1(\buffer[6][3][4] [7]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][4] [7]), .ZN(n_7_39_67));
   AOI22_X1 i_7_39_76 (.A1(\buffer[9][3][4] [7]), .A2(n_20), .B1(n_24), .B2(
      \buffer[2][3][4] [7]), .ZN(n_7_39_68));
   AOI22_X1 i_7_39_77 (.A1(\buffer[14][3][4] [7]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][4] [7]), .ZN(n_7_39_69));
   AOI22_X1 i_7_39_78 (.A1(\buffer[11][3][4] [7]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][4] [7]), .ZN(n_7_39_70));
   AOI22_X1 i_7_39_79 (.A1(\buffer[13][3][4] [7]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][3][4] [7]), .ZN(n_7_39_71));
   NAND4_X1 i_7_39_80 (.A1(n_7_39_80), .A2(n_7_39_78), .A3(n_7_39_76), .A4(
      n_7_39_72), .ZN(\output_filter[3][4] [8]));
   AOI221_X1 i_7_39_81 (.A(n_7_39_73), .B1(n_25), .B2(\buffer[0][3][4] [8]), 
      .C1(\buffer[12][3][4] [8]), .C2(n_27), .ZN(n_7_39_72));
   NAND4_X1 i_7_39_82 (.A1(n_7_39_79), .A2(n_7_39_77), .A3(n_7_39_75), .A4(
      n_7_39_74), .ZN(n_7_39_73));
   AOI22_X1 i_7_39_83 (.A1(\buffer[15][3][4] [8]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][4] [8]), .ZN(n_7_39_74));
   AOI22_X1 i_7_39_84 (.A1(\buffer[10][3][4] [8]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][4] [8]), .ZN(n_7_39_75));
   AOI22_X1 i_7_39_85 (.A1(\buffer[6][3][4] [8]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][4] [8]), .ZN(n_7_39_76));
   AOI22_X1 i_7_39_86 (.A1(\buffer[9][3][4] [8]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][3][4] [8]), .ZN(n_7_39_77));
   AOI22_X1 i_7_39_87 (.A1(\buffer[14][3][4] [8]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][4] [8]), .ZN(n_7_39_78));
   AOI22_X1 i_7_39_88 (.A1(\buffer[11][3][4] [8]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][4] [8]), .ZN(n_7_39_79));
   AOI22_X1 i_7_39_89 (.A1(\buffer[13][3][4] [8]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][4] [8]), .ZN(n_7_39_80));
   NAND4_X1 i_7_39_90 (.A1(n_7_39_89), .A2(n_7_39_87), .A3(n_7_39_85), .A4(
      n_7_39_81), .ZN(\output_filter[3][4] [9]));
   AOI221_X1 i_7_39_91 (.A(n_7_39_82), .B1(n_25), .B2(\buffer[0][3][4] [9]), 
      .C1(\buffer[12][3][4] [9]), .C2(n_27), .ZN(n_7_39_81));
   NAND4_X1 i_7_39_92 (.A1(n_7_39_88), .A2(n_7_39_86), .A3(n_7_39_84), .A4(
      n_7_39_83), .ZN(n_7_39_82));
   AOI22_X1 i_7_39_93 (.A1(\buffer[15][3][4] [9]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][4] [9]), .ZN(n_7_39_83));
   AOI22_X1 i_7_39_94 (.A1(\buffer[10][3][4] [9]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][4] [9]), .ZN(n_7_39_84));
   AOI22_X1 i_7_39_95 (.A1(\buffer[6][3][4] [9]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][4] [9]), .ZN(n_7_39_85));
   AOI22_X1 i_7_39_96 (.A1(\buffer[9][3][4] [9]), .A2(n_20), .B1(n_24), .B2(
      \buffer[2][3][4] [9]), .ZN(n_7_39_86));
   AOI22_X1 i_7_39_97 (.A1(\buffer[14][3][4] [9]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][4] [9]), .ZN(n_7_39_87));
   AOI22_X1 i_7_39_98 (.A1(\buffer[11][3][4] [9]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][4] [9]), .ZN(n_7_39_88));
   AOI22_X1 i_7_39_99 (.A1(\buffer[13][3][4] [9]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][3][4] [9]), .ZN(n_7_39_89));
   NAND4_X1 i_7_39_100 (.A1(n_7_39_98), .A2(n_7_39_96), .A3(n_7_39_94), .A4(
      n_7_39_90), .ZN(\output_filter[3][4] [10]));
   AOI221_X1 i_7_39_101 (.A(n_7_39_91), .B1(n_25), .B2(\buffer[0][3][4] [10]), 
      .C1(\buffer[12][3][4] [10]), .C2(n_27), .ZN(n_7_39_90));
   NAND4_X1 i_7_39_102 (.A1(n_7_39_97), .A2(n_7_39_95), .A3(n_7_39_93), .A4(
      n_7_39_92), .ZN(n_7_39_91));
   AOI22_X1 i_7_39_103 (.A1(\buffer[15][3][4] [10]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][4] [10]), .ZN(n_7_39_92));
   AOI22_X1 i_7_39_104 (.A1(\buffer[10][3][4] [10]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][4] [10]), .ZN(n_7_39_93));
   AOI22_X1 i_7_39_105 (.A1(\buffer[6][3][4] [10]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][4] [10]), .ZN(n_7_39_94));
   AOI22_X1 i_7_39_106 (.A1(\buffer[9][3][4] [10]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][3][4] [10]), .ZN(n_7_39_95));
   AOI22_X1 i_7_39_107 (.A1(\buffer[14][3][4] [10]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][4] [10]), .ZN(n_7_39_96));
   AOI22_X1 i_7_39_108 (.A1(\buffer[11][3][4] [10]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][4] [10]), .ZN(n_7_39_97));
   AOI22_X1 i_7_39_109 (.A1(\buffer[13][3][4] [10]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][4] [10]), .ZN(n_7_39_98));
   NAND4_X1 i_7_39_110 (.A1(n_7_39_107), .A2(n_7_39_105), .A3(n_7_39_103), 
      .A4(n_7_39_99), .ZN(\output_filter[3][4] [11]));
   AOI221_X1 i_7_39_111 (.A(n_7_39_100), .B1(n_25), .B2(\buffer[0][3][4] [11]), 
      .C1(\buffer[12][3][4] [11]), .C2(n_27), .ZN(n_7_39_99));
   NAND4_X1 i_7_39_112 (.A1(n_7_39_106), .A2(n_7_39_104), .A3(n_7_39_102), 
      .A4(n_7_39_101), .ZN(n_7_39_100));
   AOI22_X1 i_7_39_113 (.A1(\buffer[15][3][4] [11]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][4] [11]), .ZN(n_7_39_101));
   AOI22_X1 i_7_39_114 (.A1(\buffer[10][3][4] [11]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][4] [11]), .ZN(n_7_39_102));
   AOI22_X1 i_7_39_115 (.A1(\buffer[6][3][4] [11]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][4] [11]), .ZN(n_7_39_103));
   AOI22_X1 i_7_39_116 (.A1(\buffer[9][3][4] [11]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][3][4] [11]), .ZN(n_7_39_104));
   AOI22_X1 i_7_39_117 (.A1(\buffer[14][3][4] [11]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][4] [11]), .ZN(n_7_39_105));
   AOI22_X1 i_7_39_118 (.A1(\buffer[11][3][4] [11]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][4] [11]), .ZN(n_7_39_106));
   AOI22_X1 i_7_39_119 (.A1(\buffer[13][3][4] [11]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][3][4] [11]), .ZN(n_7_39_107));
   NAND4_X1 i_7_39_120 (.A1(n_7_39_116), .A2(n_7_39_114), .A3(n_7_39_112), 
      .A4(n_7_39_108), .ZN(\output_filter[3][4] [12]));
   AOI221_X1 i_7_39_121 (.A(n_7_39_109), .B1(n_25), .B2(\buffer[0][3][4] [12]), 
      .C1(\buffer[12][3][4] [12]), .C2(n_27), .ZN(n_7_39_108));
   NAND4_X1 i_7_39_122 (.A1(n_7_39_115), .A2(n_7_39_113), .A3(n_7_39_111), 
      .A4(n_7_39_110), .ZN(n_7_39_109));
   AOI22_X1 i_7_39_123 (.A1(\buffer[15][3][4] [12]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][4] [12]), .ZN(n_7_39_110));
   AOI22_X1 i_7_39_124 (.A1(\buffer[10][3][4] [12]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][4] [12]), .ZN(n_7_39_111));
   AOI22_X1 i_7_39_125 (.A1(\buffer[6][3][4] [12]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][4] [12]), .ZN(n_7_39_112));
   AOI22_X1 i_7_39_126 (.A1(\buffer[9][3][4] [12]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][3][4] [12]), .ZN(n_7_39_113));
   AOI22_X1 i_7_39_127 (.A1(\buffer[14][3][4] [12]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][4] [12]), .ZN(n_7_39_114));
   AOI22_X1 i_7_39_128 (.A1(\buffer[11][3][4] [12]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][4] [12]), .ZN(n_7_39_115));
   AOI22_X1 i_7_39_129 (.A1(\buffer[13][3][4] [12]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][4] [12]), .ZN(n_7_39_116));
   NAND4_X1 i_7_39_130 (.A1(n_7_39_125), .A2(n_7_39_123), .A3(n_7_39_121), 
      .A4(n_7_39_117), .ZN(\output_filter[3][4] [13]));
   AOI221_X1 i_7_39_131 (.A(n_7_39_118), .B1(n_25), .B2(\buffer[0][3][4] [13]), 
      .C1(\buffer[12][3][4] [13]), .C2(n_27), .ZN(n_7_39_117));
   NAND4_X1 i_7_39_132 (.A1(n_7_39_124), .A2(n_7_39_122), .A3(n_7_39_120), 
      .A4(n_7_39_119), .ZN(n_7_39_118));
   AOI22_X1 i_7_39_133 (.A1(\buffer[15][3][4] [13]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][4] [13]), .ZN(n_7_39_119));
   AOI22_X1 i_7_39_134 (.A1(\buffer[10][3][4] [13]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][4] [13]), .ZN(n_7_39_120));
   AOI22_X1 i_7_39_135 (.A1(\buffer[6][3][4] [13]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][4] [13]), .ZN(n_7_39_121));
   AOI22_X1 i_7_39_136 (.A1(\buffer[9][3][4] [13]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][3][4] [13]), .ZN(n_7_39_122));
   AOI22_X1 i_7_39_137 (.A1(\buffer[14][3][4] [13]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][4] [13]), .ZN(n_7_39_123));
   AOI22_X1 i_7_39_138 (.A1(\buffer[11][3][4] [13]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][4] [13]), .ZN(n_7_39_124));
   AOI22_X1 i_7_39_139 (.A1(\buffer[13][3][4] [13]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][3][4] [13]), .ZN(n_7_39_125));
   NAND4_X1 i_7_39_140 (.A1(n_7_39_134), .A2(n_7_39_132), .A3(n_7_39_130), 
      .A4(n_7_39_126), .ZN(\output_filter[3][4] [14]));
   AOI221_X1 i_7_39_141 (.A(n_7_39_127), .B1(n_25), .B2(\buffer[0][3][4] [14]), 
      .C1(\buffer[12][3][4] [14]), .C2(n_27), .ZN(n_7_39_126));
   NAND4_X1 i_7_39_142 (.A1(n_7_39_133), .A2(n_7_39_131), .A3(n_7_39_129), 
      .A4(n_7_39_128), .ZN(n_7_39_127));
   AOI22_X1 i_7_39_143 (.A1(\buffer[15][3][4] [14]), .A2(n_22), .B1(n_16), 
      .B2(\buffer[8][3][4] [14]), .ZN(n_7_39_128));
   AOI22_X1 i_7_39_144 (.A1(\buffer[10][3][4] [14]), .A2(n_21), .B1(n_29), 
      .B2(\buffer[7][3][4] [14]), .ZN(n_7_39_129));
   AOI22_X1 i_7_39_145 (.A1(\buffer[6][3][4] [14]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][4] [14]), .ZN(n_7_39_130));
   AOI22_X1 i_7_39_146 (.A1(\buffer[9][3][4] [14]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][3][4] [14]), .ZN(n_7_39_131));
   AOI22_X1 i_7_39_147 (.A1(\buffer[14][3][4] [14]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][4] [14]), .ZN(n_7_39_132));
   AOI22_X1 i_7_39_148 (.A1(\buffer[11][3][4] [14]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][4] [14]), .ZN(n_7_39_133));
   AOI22_X1 i_7_39_149 (.A1(\buffer[13][3][4] [14]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][4] [14]), .ZN(n_7_39_134));
   NAND2_X1 i_7_39_150 (.A1(n_7_39_137), .A2(n_7_39_135), .ZN(
      \output_filter[3][4] [15]));
   AOI221_X1 i_7_39_151 (.A(n_7_39_136), .B1(n_31), .B2(\buffer[3][3][4] [15]), 
      .C1(\buffer[14][3][4] [15]), .C2(n_19), .ZN(n_7_39_135));
   NAND3_X1 i_7_39_152 (.A1(n_7_39_143), .A2(n_7_39_141), .A3(n_7_39_139), 
      .ZN(n_7_39_136));
   AOI221_X1 i_7_39_153 (.A(n_7_39_138), .B1(n_16), .B2(\buffer[8][3][4] [15]), 
      .C1(\buffer[13][3][4] [15]), .C2(n_26), .ZN(n_7_39_137));
   NAND3_X1 i_7_39_154 (.A1(n_7_39_144), .A2(n_7_39_142), .A3(n_7_39_140), 
      .ZN(n_7_39_138));
   AOI22_X1 i_7_39_155 (.A1(\buffer[11][3][4] [15]), .A2(n_17), .B1(n_24), 
      .B2(\buffer[2][3][4] [15]), .ZN(n_7_39_139));
   AOI22_X1 i_7_39_156 (.A1(\buffer[10][3][4] [15]), .A2(n_21), .B1(n_23), 
      .B2(\buffer[1][3][4] [15]), .ZN(n_7_39_140));
   AOI22_X1 i_7_39_157 (.A1(\buffer[6][3][4] [15]), .A2(n_28), .B1(n_18), 
      .B2(\buffer[5][3][4] [15]), .ZN(n_7_39_141));
   AOI22_X1 i_7_39_158 (.A1(\buffer[9][3][4] [15]), .A2(n_20), .B1(n_30), 
      .B2(\buffer[4][3][4] [15]), .ZN(n_7_39_142));
   AOI22_X1 i_7_39_159 (.A1(\buffer[7][3][4] [15]), .A2(n_29), .B1(n_25), 
      .B2(\buffer[0][3][4] [15]), .ZN(n_7_39_143));
   AOI22_X1 i_7_39_160 (.A1(\buffer[15][3][4] [15]), .A2(n_22), .B1(n_27), 
      .B2(\buffer[12][3][4] [15]), .ZN(n_7_39_144));
   NAND4_X1 i_8_37_0 (.A1(n_8_37_8), .A2(n_8_37_6), .A3(n_8_37_4), .A4(n_8_37_0), 
      .ZN(\output_filter[3][2] [0]));
   AOI221_X1 i_8_37_1 (.A(n_8_37_1), .B1(n_25), .B2(\buffer[0][3][2] [0]), 
      .C1(\buffer[12][3][2] [0]), .C2(n_27), .ZN(n_8_37_0));
   NAND4_X1 i_8_37_2 (.A1(n_8_37_7), .A2(n_8_37_5), .A3(n_8_37_3), .A4(n_8_37_2), 
      .ZN(n_8_37_1));
   AOI22_X1 i_8_37_3 (.A1(\buffer[15][3][2] [0]), .A2(n_22), .B1(n_29), .B2(
      \buffer[7][3][2] [0]), .ZN(n_8_37_2));
   AOI22_X1 i_8_37_4 (.A1(\buffer[10][3][2] [0]), .A2(n_21), .B1(n_16), .B2(
      \buffer[8][3][2] [0]), .ZN(n_8_37_3));
   AOI22_X1 i_8_37_5 (.A1(\buffer[6][3][2] [0]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][2] [0]), .ZN(n_8_37_4));
   AOI22_X1 i_8_37_6 (.A1(\buffer[9][3][2] [0]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][3][2] [0]), .ZN(n_8_37_5));
   AOI22_X1 i_8_37_7 (.A1(\buffer[14][3][2] [0]), .A2(n_19), .B1(n_23), .B2(
      \buffer[1][3][2] [0]), .ZN(n_8_37_6));
   AOI22_X1 i_8_37_8 (.A1(\buffer[11][3][2] [0]), .A2(n_17), .B1(n_18), .B2(
      \buffer[5][3][2] [0]), .ZN(n_8_37_7));
   AOI22_X1 i_8_37_9 (.A1(\buffer[13][3][2] [0]), .A2(n_26), .B1(n_24), .B2(
      \buffer[2][3][2] [0]), .ZN(n_8_37_8));
   NAND4_X1 i_8_37_10 (.A1(n_8_37_17), .A2(n_8_37_15), .A3(n_8_37_13), .A4(
      n_8_37_9), .ZN(\output_filter[3][2] [1]));
   AOI221_X1 i_8_37_11 (.A(n_8_37_10), .B1(n_25), .B2(\buffer[0][3][2] [1]), 
      .C1(\buffer[12][3][2] [1]), .C2(n_27), .ZN(n_8_37_9));
   NAND4_X1 i_8_37_12 (.A1(n_8_37_16), .A2(n_8_37_14), .A3(n_8_37_12), .A4(
      n_8_37_11), .ZN(n_8_37_10));
   AOI22_X1 i_8_37_13 (.A1(\buffer[15][3][2] [1]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][2] [1]), .ZN(n_8_37_11));
   AOI22_X1 i_8_37_14 (.A1(\buffer[10][3][2] [1]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][2] [1]), .ZN(n_8_37_12));
   AOI22_X1 i_8_37_15 (.A1(\buffer[6][3][2] [1]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][2] [1]), .ZN(n_8_37_13));
   AOI22_X1 i_8_37_16 (.A1(\buffer[9][3][2] [1]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][3][2] [1]), .ZN(n_8_37_14));
   AOI22_X1 i_8_37_17 (.A1(\buffer[14][3][2] [1]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][2] [1]), .ZN(n_8_37_15));
   AOI22_X1 i_8_37_18 (.A1(\buffer[11][3][2] [1]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][2] [1]), .ZN(n_8_37_16));
   AOI22_X1 i_8_37_19 (.A1(\buffer[13][3][2] [1]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][2] [1]), .ZN(n_8_37_17));
   NAND4_X1 i_8_37_20 (.A1(n_8_37_26), .A2(n_8_37_24), .A3(n_8_37_22), .A4(
      n_8_37_18), .ZN(\output_filter[3][2] [2]));
   AOI221_X1 i_8_37_21 (.A(n_8_37_19), .B1(n_25), .B2(\buffer[0][3][2] [2]), 
      .C1(\buffer[12][3][2] [2]), .C2(n_27), .ZN(n_8_37_18));
   NAND4_X1 i_8_37_22 (.A1(n_8_37_25), .A2(n_8_37_23), .A3(n_8_37_21), .A4(
      n_8_37_20), .ZN(n_8_37_19));
   AOI22_X1 i_8_37_23 (.A1(\buffer[15][3][2] [2]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][2] [2]), .ZN(n_8_37_20));
   AOI22_X1 i_8_37_24 (.A1(\buffer[10][3][2] [2]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][2] [2]), .ZN(n_8_37_21));
   AOI22_X1 i_8_37_25 (.A1(\buffer[6][3][2] [2]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][2] [2]), .ZN(n_8_37_22));
   AOI22_X1 i_8_37_26 (.A1(\buffer[9][3][2] [2]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][3][2] [2]), .ZN(n_8_37_23));
   AOI22_X1 i_8_37_27 (.A1(\buffer[14][3][2] [2]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][2] [2]), .ZN(n_8_37_24));
   AOI22_X1 i_8_37_28 (.A1(\buffer[11][3][2] [2]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][2] [2]), .ZN(n_8_37_25));
   AOI22_X1 i_8_37_29 (.A1(\buffer[13][3][2] [2]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][2] [2]), .ZN(n_8_37_26));
   NAND4_X1 i_8_37_30 (.A1(n_8_37_35), .A2(n_8_37_33), .A3(n_8_37_31), .A4(
      n_8_37_27), .ZN(\output_filter[3][2] [3]));
   AOI221_X1 i_8_37_31 (.A(n_8_37_28), .B1(n_25), .B2(\buffer[0][3][2] [3]), 
      .C1(\buffer[12][3][2] [3]), .C2(n_27), .ZN(n_8_37_27));
   NAND4_X1 i_8_37_32 (.A1(n_8_37_34), .A2(n_8_37_32), .A3(n_8_37_30), .A4(
      n_8_37_29), .ZN(n_8_37_28));
   AOI22_X1 i_8_37_33 (.A1(\buffer[15][3][2] [3]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][2] [3]), .ZN(n_8_37_29));
   AOI22_X1 i_8_37_34 (.A1(\buffer[10][3][2] [3]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][2] [3]), .ZN(n_8_37_30));
   AOI22_X1 i_8_37_35 (.A1(\buffer[6][3][2] [3]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][2] [3]), .ZN(n_8_37_31));
   AOI22_X1 i_8_37_36 (.A1(\buffer[9][3][2] [3]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][3][2] [3]), .ZN(n_8_37_32));
   AOI22_X1 i_8_37_37 (.A1(\buffer[14][3][2] [3]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][2] [3]), .ZN(n_8_37_33));
   AOI22_X1 i_8_37_38 (.A1(\buffer[11][3][2] [3]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][2] [3]), .ZN(n_8_37_34));
   AOI22_X1 i_8_37_39 (.A1(\buffer[13][3][2] [3]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][2] [3]), .ZN(n_8_37_35));
   NAND4_X1 i_8_37_40 (.A1(n_8_37_44), .A2(n_8_37_42), .A3(n_8_37_40), .A4(
      n_8_37_36), .ZN(\output_filter[3][2] [4]));
   AOI221_X1 i_8_37_41 (.A(n_8_37_37), .B1(n_25), .B2(\buffer[0][3][2] [4]), 
      .C1(\buffer[12][3][2] [4]), .C2(n_27), .ZN(n_8_37_36));
   NAND4_X1 i_8_37_42 (.A1(n_8_37_43), .A2(n_8_37_41), .A3(n_8_37_39), .A4(
      n_8_37_38), .ZN(n_8_37_37));
   AOI22_X1 i_8_37_43 (.A1(\buffer[15][3][2] [4]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][2] [4]), .ZN(n_8_37_38));
   AOI22_X1 i_8_37_44 (.A1(\buffer[10][3][2] [4]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][2] [4]), .ZN(n_8_37_39));
   AOI22_X1 i_8_37_45 (.A1(\buffer[6][3][2] [4]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][2] [4]), .ZN(n_8_37_40));
   AOI22_X1 i_8_37_46 (.A1(\buffer[9][3][2] [4]), .A2(n_20), .B1(n_24), .B2(
      \buffer[2][3][2] [4]), .ZN(n_8_37_41));
   AOI22_X1 i_8_37_47 (.A1(\buffer[14][3][2] [4]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][2] [4]), .ZN(n_8_37_42));
   AOI22_X1 i_8_37_48 (.A1(\buffer[11][3][2] [4]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][2] [4]), .ZN(n_8_37_43));
   AOI22_X1 i_8_37_49 (.A1(\buffer[13][3][2] [4]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][3][2] [4]), .ZN(n_8_37_44));
   NAND4_X1 i_8_37_50 (.A1(n_8_37_53), .A2(n_8_37_51), .A3(n_8_37_49), .A4(
      n_8_37_45), .ZN(\output_filter[3][2] [5]));
   AOI221_X1 i_8_37_51 (.A(n_8_37_46), .B1(n_25), .B2(\buffer[0][3][2] [5]), 
      .C1(\buffer[12][3][2] [5]), .C2(n_27), .ZN(n_8_37_45));
   NAND4_X1 i_8_37_52 (.A1(n_8_37_52), .A2(n_8_37_50), .A3(n_8_37_48), .A4(
      n_8_37_47), .ZN(n_8_37_46));
   AOI22_X1 i_8_37_53 (.A1(\buffer[15][3][2] [5]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][2] [5]), .ZN(n_8_37_47));
   AOI22_X1 i_8_37_54 (.A1(\buffer[10][3][2] [5]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][2] [5]), .ZN(n_8_37_48));
   AOI22_X1 i_8_37_55 (.A1(\buffer[6][3][2] [5]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][2] [5]), .ZN(n_8_37_49));
   AOI22_X1 i_8_37_56 (.A1(\buffer[9][3][2] [5]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][3][2] [5]), .ZN(n_8_37_50));
   AOI22_X1 i_8_37_57 (.A1(\buffer[14][3][2] [5]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][2] [5]), .ZN(n_8_37_51));
   AOI22_X1 i_8_37_58 (.A1(\buffer[11][3][2] [5]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][2] [5]), .ZN(n_8_37_52));
   AOI22_X1 i_8_37_59 (.A1(\buffer[13][3][2] [5]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][2] [5]), .ZN(n_8_37_53));
   NAND4_X1 i_8_37_60 (.A1(n_8_37_62), .A2(n_8_37_60), .A3(n_8_37_58), .A4(
      n_8_37_54), .ZN(\output_filter[3][2] [6]));
   AOI221_X1 i_8_37_61 (.A(n_8_37_55), .B1(n_25), .B2(\buffer[0][3][2] [6]), 
      .C1(\buffer[12][3][2] [6]), .C2(n_27), .ZN(n_8_37_54));
   NAND4_X1 i_8_37_62 (.A1(n_8_37_61), .A2(n_8_37_59), .A3(n_8_37_57), .A4(
      n_8_37_56), .ZN(n_8_37_55));
   AOI22_X1 i_8_37_63 (.A1(\buffer[15][3][2] [6]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][2] [6]), .ZN(n_8_37_56));
   AOI22_X1 i_8_37_64 (.A1(\buffer[10][3][2] [6]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][2] [6]), .ZN(n_8_37_57));
   AOI22_X1 i_8_37_65 (.A1(\buffer[6][3][2] [6]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][2] [6]), .ZN(n_8_37_58));
   AOI22_X1 i_8_37_66 (.A1(\buffer[9][3][2] [6]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][3][2] [6]), .ZN(n_8_37_59));
   AOI22_X1 i_8_37_67 (.A1(\buffer[14][3][2] [6]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][2] [6]), .ZN(n_8_37_60));
   AOI22_X1 i_8_37_68 (.A1(\buffer[11][3][2] [6]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][2] [6]), .ZN(n_8_37_61));
   AOI22_X1 i_8_37_69 (.A1(\buffer[13][3][2] [6]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][2] [6]), .ZN(n_8_37_62));
   NAND4_X1 i_8_37_70 (.A1(n_8_37_71), .A2(n_8_37_69), .A3(n_8_37_67), .A4(
      n_8_37_63), .ZN(\output_filter[3][2] [7]));
   AOI221_X1 i_8_37_71 (.A(n_8_37_64), .B1(n_25), .B2(\buffer[0][3][2] [7]), 
      .C1(\buffer[12][3][2] [7]), .C2(n_27), .ZN(n_8_37_63));
   NAND4_X1 i_8_37_72 (.A1(n_8_37_70), .A2(n_8_37_68), .A3(n_8_37_66), .A4(
      n_8_37_65), .ZN(n_8_37_64));
   AOI22_X1 i_8_37_73 (.A1(\buffer[15][3][2] [7]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][2] [7]), .ZN(n_8_37_65));
   AOI22_X1 i_8_37_74 (.A1(\buffer[10][3][2] [7]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][2] [7]), .ZN(n_8_37_66));
   AOI22_X1 i_8_37_75 (.A1(\buffer[6][3][2] [7]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][2] [7]), .ZN(n_8_37_67));
   AOI22_X1 i_8_37_76 (.A1(\buffer[9][3][2] [7]), .A2(n_20), .B1(n_24), .B2(
      \buffer[2][3][2] [7]), .ZN(n_8_37_68));
   AOI22_X1 i_8_37_77 (.A1(\buffer[14][3][2] [7]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][2] [7]), .ZN(n_8_37_69));
   AOI22_X1 i_8_37_78 (.A1(\buffer[11][3][2] [7]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][2] [7]), .ZN(n_8_37_70));
   AOI22_X1 i_8_37_79 (.A1(\buffer[13][3][2] [7]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][3][2] [7]), .ZN(n_8_37_71));
   NAND4_X1 i_8_37_80 (.A1(n_8_37_80), .A2(n_8_37_78), .A3(n_8_37_76), .A4(
      n_8_37_72), .ZN(\output_filter[3][2] [8]));
   AOI221_X1 i_8_37_81 (.A(n_8_37_73), .B1(n_25), .B2(\buffer[0][3][2] [8]), 
      .C1(\buffer[12][3][2] [8]), .C2(n_27), .ZN(n_8_37_72));
   NAND4_X1 i_8_37_82 (.A1(n_8_37_79), .A2(n_8_37_77), .A3(n_8_37_75), .A4(
      n_8_37_74), .ZN(n_8_37_73));
   AOI22_X1 i_8_37_83 (.A1(\buffer[15][3][2] [8]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][2] [8]), .ZN(n_8_37_74));
   AOI22_X1 i_8_37_84 (.A1(\buffer[10][3][2] [8]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][2] [8]), .ZN(n_8_37_75));
   AOI22_X1 i_8_37_85 (.A1(\buffer[6][3][2] [8]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][2] [8]), .ZN(n_8_37_76));
   AOI22_X1 i_8_37_86 (.A1(\buffer[9][3][2] [8]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][3][2] [8]), .ZN(n_8_37_77));
   AOI22_X1 i_8_37_87 (.A1(\buffer[14][3][2] [8]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][2] [8]), .ZN(n_8_37_78));
   AOI22_X1 i_8_37_88 (.A1(\buffer[11][3][2] [8]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][2] [8]), .ZN(n_8_37_79));
   AOI22_X1 i_8_37_89 (.A1(\buffer[13][3][2] [8]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][2] [8]), .ZN(n_8_37_80));
   NAND4_X1 i_8_37_90 (.A1(n_8_37_89), .A2(n_8_37_87), .A3(n_8_37_85), .A4(
      n_8_37_81), .ZN(\output_filter[3][2] [9]));
   AOI221_X1 i_8_37_91 (.A(n_8_37_82), .B1(n_25), .B2(\buffer[0][3][2] [9]), 
      .C1(\buffer[12][3][2] [9]), .C2(n_27), .ZN(n_8_37_81));
   NAND4_X1 i_8_37_92 (.A1(n_8_37_88), .A2(n_8_37_86), .A3(n_8_37_84), .A4(
      n_8_37_83), .ZN(n_8_37_82));
   AOI22_X1 i_8_37_93 (.A1(\buffer[15][3][2] [9]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][2] [9]), .ZN(n_8_37_83));
   AOI22_X1 i_8_37_94 (.A1(\buffer[10][3][2] [9]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][2] [9]), .ZN(n_8_37_84));
   AOI22_X1 i_8_37_95 (.A1(\buffer[6][3][2] [9]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][2] [9]), .ZN(n_8_37_85));
   AOI22_X1 i_8_37_96 (.A1(\buffer[9][3][2] [9]), .A2(n_20), .B1(n_24), .B2(
      \buffer[2][3][2] [9]), .ZN(n_8_37_86));
   AOI22_X1 i_8_37_97 (.A1(\buffer[14][3][2] [9]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][2] [9]), .ZN(n_8_37_87));
   AOI22_X1 i_8_37_98 (.A1(\buffer[11][3][2] [9]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][2] [9]), .ZN(n_8_37_88));
   AOI22_X1 i_8_37_99 (.A1(\buffer[13][3][2] [9]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][3][2] [9]), .ZN(n_8_37_89));
   NAND4_X1 i_8_37_100 (.A1(n_8_37_98), .A2(n_8_37_96), .A3(n_8_37_94), .A4(
      n_8_37_90), .ZN(\output_filter[3][2] [10]));
   AOI221_X1 i_8_37_101 (.A(n_8_37_91), .B1(n_25), .B2(\buffer[0][3][2] [10]), 
      .C1(\buffer[12][3][2] [10]), .C2(n_27), .ZN(n_8_37_90));
   NAND4_X1 i_8_37_102 (.A1(n_8_37_97), .A2(n_8_37_95), .A3(n_8_37_93), .A4(
      n_8_37_92), .ZN(n_8_37_91));
   AOI22_X1 i_8_37_103 (.A1(\buffer[15][3][2] [10]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][2] [10]), .ZN(n_8_37_92));
   AOI22_X1 i_8_37_104 (.A1(\buffer[10][3][2] [10]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][2] [10]), .ZN(n_8_37_93));
   AOI22_X1 i_8_37_105 (.A1(\buffer[6][3][2] [10]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][2] [10]), .ZN(n_8_37_94));
   AOI22_X1 i_8_37_106 (.A1(\buffer[9][3][2] [10]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][3][2] [10]), .ZN(n_8_37_95));
   AOI22_X1 i_8_37_107 (.A1(\buffer[14][3][2] [10]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][2] [10]), .ZN(n_8_37_96));
   AOI22_X1 i_8_37_108 (.A1(\buffer[11][3][2] [10]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][2] [10]), .ZN(n_8_37_97));
   AOI22_X1 i_8_37_109 (.A1(\buffer[13][3][2] [10]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][2] [10]), .ZN(n_8_37_98));
   NAND4_X1 i_8_37_110 (.A1(n_8_37_107), .A2(n_8_37_105), .A3(n_8_37_103), 
      .A4(n_8_37_99), .ZN(\output_filter[3][2] [11]));
   AOI221_X1 i_8_37_111 (.A(n_8_37_100), .B1(n_25), .B2(\buffer[0][3][2] [11]), 
      .C1(\buffer[12][3][2] [11]), .C2(n_27), .ZN(n_8_37_99));
   NAND4_X1 i_8_37_112 (.A1(n_8_37_106), .A2(n_8_37_104), .A3(n_8_37_102), 
      .A4(n_8_37_101), .ZN(n_8_37_100));
   AOI22_X1 i_8_37_113 (.A1(\buffer[15][3][2] [11]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][2] [11]), .ZN(n_8_37_101));
   AOI22_X1 i_8_37_114 (.A1(\buffer[10][3][2] [11]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][2] [11]), .ZN(n_8_37_102));
   AOI22_X1 i_8_37_115 (.A1(\buffer[6][3][2] [11]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][2] [11]), .ZN(n_8_37_103));
   AOI22_X1 i_8_37_116 (.A1(\buffer[9][3][2] [11]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][3][2] [11]), .ZN(n_8_37_104));
   AOI22_X1 i_8_37_117 (.A1(\buffer[14][3][2] [11]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][2] [11]), .ZN(n_8_37_105));
   AOI22_X1 i_8_37_118 (.A1(\buffer[11][3][2] [11]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][2] [11]), .ZN(n_8_37_106));
   AOI22_X1 i_8_37_119 (.A1(\buffer[13][3][2] [11]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][3][2] [11]), .ZN(n_8_37_107));
   NAND4_X1 i_8_37_120 (.A1(n_8_37_116), .A2(n_8_37_114), .A3(n_8_37_112), 
      .A4(n_8_37_108), .ZN(\output_filter[3][2] [12]));
   AOI221_X1 i_8_37_121 (.A(n_8_37_109), .B1(n_25), .B2(\buffer[0][3][2] [12]), 
      .C1(\buffer[12][3][2] [12]), .C2(n_27), .ZN(n_8_37_108));
   NAND4_X1 i_8_37_122 (.A1(n_8_37_115), .A2(n_8_37_113), .A3(n_8_37_111), 
      .A4(n_8_37_110), .ZN(n_8_37_109));
   AOI22_X1 i_8_37_123 (.A1(\buffer[15][3][2] [12]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][2] [12]), .ZN(n_8_37_110));
   AOI22_X1 i_8_37_124 (.A1(\buffer[10][3][2] [12]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][2] [12]), .ZN(n_8_37_111));
   AOI22_X1 i_8_37_125 (.A1(\buffer[6][3][2] [12]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][2] [12]), .ZN(n_8_37_112));
   AOI22_X1 i_8_37_126 (.A1(\buffer[9][3][2] [12]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][3][2] [12]), .ZN(n_8_37_113));
   AOI22_X1 i_8_37_127 (.A1(\buffer[14][3][2] [12]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][2] [12]), .ZN(n_8_37_114));
   AOI22_X1 i_8_37_128 (.A1(\buffer[11][3][2] [12]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][2] [12]), .ZN(n_8_37_115));
   AOI22_X1 i_8_37_129 (.A1(\buffer[13][3][2] [12]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][2] [12]), .ZN(n_8_37_116));
   NAND4_X1 i_8_37_130 (.A1(n_8_37_125), .A2(n_8_37_123), .A3(n_8_37_121), 
      .A4(n_8_37_117), .ZN(\output_filter[3][2] [13]));
   AOI221_X1 i_8_37_131 (.A(n_8_37_118), .B1(n_25), .B2(\buffer[0][3][2] [13]), 
      .C1(\buffer[12][3][2] [13]), .C2(n_27), .ZN(n_8_37_117));
   NAND4_X1 i_8_37_132 (.A1(n_8_37_124), .A2(n_8_37_122), .A3(n_8_37_120), 
      .A4(n_8_37_119), .ZN(n_8_37_118));
   AOI22_X1 i_8_37_133 (.A1(\buffer[15][3][2] [13]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][2] [13]), .ZN(n_8_37_119));
   AOI22_X1 i_8_37_134 (.A1(\buffer[10][3][2] [13]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][2] [13]), .ZN(n_8_37_120));
   AOI22_X1 i_8_37_135 (.A1(\buffer[6][3][2] [13]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][2] [13]), .ZN(n_8_37_121));
   AOI22_X1 i_8_37_136 (.A1(\buffer[9][3][2] [13]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][3][2] [13]), .ZN(n_8_37_122));
   AOI22_X1 i_8_37_137 (.A1(\buffer[14][3][2] [13]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][2] [13]), .ZN(n_8_37_123));
   AOI22_X1 i_8_37_138 (.A1(\buffer[11][3][2] [13]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][2] [13]), .ZN(n_8_37_124));
   AOI22_X1 i_8_37_139 (.A1(\buffer[13][3][2] [13]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][3][2] [13]), .ZN(n_8_37_125));
   NAND4_X1 i_8_37_140 (.A1(n_8_37_134), .A2(n_8_37_132), .A3(n_8_37_130), 
      .A4(n_8_37_126), .ZN(\output_filter[3][2] [14]));
   AOI221_X1 i_8_37_141 (.A(n_8_37_127), .B1(n_25), .B2(\buffer[0][3][2] [14]), 
      .C1(\buffer[12][3][2] [14]), .C2(n_27), .ZN(n_8_37_126));
   NAND4_X1 i_8_37_142 (.A1(n_8_37_133), .A2(n_8_37_131), .A3(n_8_37_129), 
      .A4(n_8_37_128), .ZN(n_8_37_127));
   AOI22_X1 i_8_37_143 (.A1(\buffer[15][3][2] [14]), .A2(n_22), .B1(n_16), 
      .B2(\buffer[8][3][2] [14]), .ZN(n_8_37_128));
   AOI22_X1 i_8_37_144 (.A1(\buffer[10][3][2] [14]), .A2(n_21), .B1(n_29), 
      .B2(\buffer[7][3][2] [14]), .ZN(n_8_37_129));
   AOI22_X1 i_8_37_145 (.A1(\buffer[6][3][2] [14]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][2] [14]), .ZN(n_8_37_130));
   AOI22_X1 i_8_37_146 (.A1(\buffer[9][3][2] [14]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][3][2] [14]), .ZN(n_8_37_131));
   AOI22_X1 i_8_37_147 (.A1(\buffer[14][3][2] [14]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][2] [14]), .ZN(n_8_37_132));
   AOI22_X1 i_8_37_148 (.A1(\buffer[11][3][2] [14]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][2] [14]), .ZN(n_8_37_133));
   AOI22_X1 i_8_37_149 (.A1(\buffer[13][3][2] [14]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][2] [14]), .ZN(n_8_37_134));
   NAND2_X1 i_8_37_150 (.A1(n_8_37_137), .A2(n_8_37_135), .ZN(
      \output_filter[3][2] [15]));
   AOI221_X1 i_8_37_151 (.A(n_8_37_136), .B1(n_31), .B2(\buffer[3][3][2] [15]), 
      .C1(\buffer[14][3][2] [15]), .C2(n_19), .ZN(n_8_37_135));
   NAND3_X1 i_8_37_152 (.A1(n_8_37_143), .A2(n_8_37_141), .A3(n_8_37_139), 
      .ZN(n_8_37_136));
   AOI221_X1 i_8_37_153 (.A(n_8_37_138), .B1(n_16), .B2(\buffer[8][3][2] [15]), 
      .C1(\buffer[13][3][2] [15]), .C2(n_26), .ZN(n_8_37_137));
   NAND3_X1 i_8_37_154 (.A1(n_8_37_144), .A2(n_8_37_142), .A3(n_8_37_140), 
      .ZN(n_8_37_138));
   AOI22_X1 i_8_37_155 (.A1(\buffer[11][3][2] [15]), .A2(n_17), .B1(n_24), 
      .B2(\buffer[2][3][2] [15]), .ZN(n_8_37_139));
   AOI22_X1 i_8_37_156 (.A1(\buffer[10][3][2] [15]), .A2(n_21), .B1(n_23), 
      .B2(\buffer[1][3][2] [15]), .ZN(n_8_37_140));
   AOI22_X1 i_8_37_157 (.A1(\buffer[6][3][2] [15]), .A2(n_28), .B1(n_18), 
      .B2(\buffer[5][3][2] [15]), .ZN(n_8_37_141));
   AOI22_X1 i_8_37_158 (.A1(\buffer[9][3][2] [15]), .A2(n_20), .B1(n_30), 
      .B2(\buffer[4][3][2] [15]), .ZN(n_8_37_142));
   AOI22_X1 i_8_37_159 (.A1(\buffer[7][3][2] [15]), .A2(n_29), .B1(n_25), 
      .B2(\buffer[0][3][2] [15]), .ZN(n_8_37_143));
   AOI22_X1 i_8_37_160 (.A1(\buffer[15][3][2] [15]), .A2(n_22), .B1(n_27), 
      .B2(\buffer[12][3][2] [15]), .ZN(n_8_37_144));
   NAND4_X1 i_9_36_0 (.A1(n_9_36_8), .A2(n_9_36_6), .A3(n_9_36_4), .A4(n_9_36_0), 
      .ZN(\output_filter[3][1] [0]));
   AOI221_X1 i_9_36_1 (.A(n_9_36_1), .B1(n_25), .B2(\buffer[0][3][1] [0]), 
      .C1(\buffer[12][3][1] [0]), .C2(n_27), .ZN(n_9_36_0));
   NAND4_X1 i_9_36_2 (.A1(n_9_36_7), .A2(n_9_36_5), .A3(n_9_36_3), .A4(n_9_36_2), 
      .ZN(n_9_36_1));
   AOI22_X1 i_9_36_3 (.A1(\buffer[15][3][1] [0]), .A2(n_22), .B1(n_29), .B2(
      \buffer[7][3][1] [0]), .ZN(n_9_36_2));
   AOI22_X1 i_9_36_4 (.A1(\buffer[10][3][1] [0]), .A2(n_21), .B1(n_16), .B2(
      \buffer[8][3][1] [0]), .ZN(n_9_36_3));
   AOI22_X1 i_9_36_5 (.A1(\buffer[6][3][1] [0]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][1] [0]), .ZN(n_9_36_4));
   AOI22_X1 i_9_36_6 (.A1(\buffer[9][3][1] [0]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][3][1] [0]), .ZN(n_9_36_5));
   AOI22_X1 i_9_36_7 (.A1(\buffer[14][3][1] [0]), .A2(n_19), .B1(n_23), .B2(
      \buffer[1][3][1] [0]), .ZN(n_9_36_6));
   AOI22_X1 i_9_36_8 (.A1(\buffer[11][3][1] [0]), .A2(n_17), .B1(n_18), .B2(
      \buffer[5][3][1] [0]), .ZN(n_9_36_7));
   AOI22_X1 i_9_36_9 (.A1(\buffer[13][3][1] [0]), .A2(n_26), .B1(n_24), .B2(
      \buffer[2][3][1] [0]), .ZN(n_9_36_8));
   NAND4_X1 i_9_36_10 (.A1(n_9_36_17), .A2(n_9_36_15), .A3(n_9_36_13), .A4(
      n_9_36_9), .ZN(\output_filter[3][1] [1]));
   AOI221_X1 i_9_36_11 (.A(n_9_36_10), .B1(n_25), .B2(\buffer[0][3][1] [1]), 
      .C1(\buffer[12][3][1] [1]), .C2(n_27), .ZN(n_9_36_9));
   NAND4_X1 i_9_36_12 (.A1(n_9_36_16), .A2(n_9_36_14), .A3(n_9_36_12), .A4(
      n_9_36_11), .ZN(n_9_36_10));
   AOI22_X1 i_9_36_13 (.A1(\buffer[15][3][1] [1]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][1] [1]), .ZN(n_9_36_11));
   AOI22_X1 i_9_36_14 (.A1(\buffer[10][3][1] [1]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][1] [1]), .ZN(n_9_36_12));
   AOI22_X1 i_9_36_15 (.A1(\buffer[6][3][1] [1]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][1] [1]), .ZN(n_9_36_13));
   AOI22_X1 i_9_36_16 (.A1(\buffer[9][3][1] [1]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][3][1] [1]), .ZN(n_9_36_14));
   AOI22_X1 i_9_36_17 (.A1(\buffer[14][3][1] [1]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][1] [1]), .ZN(n_9_36_15));
   AOI22_X1 i_9_36_18 (.A1(\buffer[11][3][1] [1]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][1] [1]), .ZN(n_9_36_16));
   AOI22_X1 i_9_36_19 (.A1(\buffer[13][3][1] [1]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][1] [1]), .ZN(n_9_36_17));
   NAND4_X1 i_9_36_20 (.A1(n_9_36_26), .A2(n_9_36_24), .A3(n_9_36_22), .A4(
      n_9_36_18), .ZN(\output_filter[3][1] [2]));
   AOI221_X1 i_9_36_21 (.A(n_9_36_19), .B1(n_25), .B2(\buffer[0][3][1] [2]), 
      .C1(\buffer[12][3][1] [2]), .C2(n_27), .ZN(n_9_36_18));
   NAND4_X1 i_9_36_22 (.A1(n_9_36_25), .A2(n_9_36_23), .A3(n_9_36_21), .A4(
      n_9_36_20), .ZN(n_9_36_19));
   AOI22_X1 i_9_36_23 (.A1(\buffer[15][3][1] [2]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][1] [2]), .ZN(n_9_36_20));
   AOI22_X1 i_9_36_24 (.A1(\buffer[10][3][1] [2]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][1] [2]), .ZN(n_9_36_21));
   AOI22_X1 i_9_36_25 (.A1(\buffer[6][3][1] [2]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][1] [2]), .ZN(n_9_36_22));
   AOI22_X1 i_9_36_26 (.A1(\buffer[9][3][1] [2]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][3][1] [2]), .ZN(n_9_36_23));
   AOI22_X1 i_9_36_27 (.A1(\buffer[14][3][1] [2]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][1] [2]), .ZN(n_9_36_24));
   AOI22_X1 i_9_36_28 (.A1(\buffer[11][3][1] [2]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][1] [2]), .ZN(n_9_36_25));
   AOI22_X1 i_9_36_29 (.A1(\buffer[13][3][1] [2]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][1] [2]), .ZN(n_9_36_26));
   NAND4_X1 i_9_36_30 (.A1(n_9_36_35), .A2(n_9_36_33), .A3(n_9_36_31), .A4(
      n_9_36_27), .ZN(\output_filter[3][1] [3]));
   AOI221_X1 i_9_36_31 (.A(n_9_36_28), .B1(n_25), .B2(\buffer[0][3][1] [3]), 
      .C1(\buffer[12][3][1] [3]), .C2(n_27), .ZN(n_9_36_27));
   NAND4_X1 i_9_36_32 (.A1(n_9_36_34), .A2(n_9_36_32), .A3(n_9_36_30), .A4(
      n_9_36_29), .ZN(n_9_36_28));
   AOI22_X1 i_9_36_33 (.A1(\buffer[15][3][1] [3]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][1] [3]), .ZN(n_9_36_29));
   AOI22_X1 i_9_36_34 (.A1(\buffer[10][3][1] [3]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][1] [3]), .ZN(n_9_36_30));
   AOI22_X1 i_9_36_35 (.A1(\buffer[6][3][1] [3]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][1] [3]), .ZN(n_9_36_31));
   AOI22_X1 i_9_36_36 (.A1(\buffer[9][3][1] [3]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][3][1] [3]), .ZN(n_9_36_32));
   AOI22_X1 i_9_36_37 (.A1(\buffer[14][3][1] [3]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][1] [3]), .ZN(n_9_36_33));
   AOI22_X1 i_9_36_38 (.A1(\buffer[11][3][1] [3]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][1] [3]), .ZN(n_9_36_34));
   AOI22_X1 i_9_36_39 (.A1(\buffer[13][3][1] [3]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][1] [3]), .ZN(n_9_36_35));
   NAND4_X1 i_9_36_40 (.A1(n_9_36_44), .A2(n_9_36_42), .A3(n_9_36_40), .A4(
      n_9_36_36), .ZN(\output_filter[3][1] [4]));
   AOI221_X1 i_9_36_41 (.A(n_9_36_37), .B1(n_25), .B2(\buffer[0][3][1] [4]), 
      .C1(\buffer[12][3][1] [4]), .C2(n_27), .ZN(n_9_36_36));
   NAND4_X1 i_9_36_42 (.A1(n_9_36_43), .A2(n_9_36_41), .A3(n_9_36_39), .A4(
      n_9_36_38), .ZN(n_9_36_37));
   AOI22_X1 i_9_36_43 (.A1(\buffer[15][3][1] [4]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][1] [4]), .ZN(n_9_36_38));
   AOI22_X1 i_9_36_44 (.A1(\buffer[10][3][1] [4]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][1] [4]), .ZN(n_9_36_39));
   AOI22_X1 i_9_36_45 (.A1(\buffer[6][3][1] [4]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][1] [4]), .ZN(n_9_36_40));
   AOI22_X1 i_9_36_46 (.A1(\buffer[9][3][1] [4]), .A2(n_20), .B1(n_24), .B2(
      \buffer[2][3][1] [4]), .ZN(n_9_36_41));
   AOI22_X1 i_9_36_47 (.A1(\buffer[14][3][1] [4]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][1] [4]), .ZN(n_9_36_42));
   AOI22_X1 i_9_36_48 (.A1(\buffer[11][3][1] [4]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][1] [4]), .ZN(n_9_36_43));
   AOI22_X1 i_9_36_49 (.A1(\buffer[13][3][1] [4]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][3][1] [4]), .ZN(n_9_36_44));
   NAND4_X1 i_9_36_50 (.A1(n_9_36_53), .A2(n_9_36_51), .A3(n_9_36_49), .A4(
      n_9_36_45), .ZN(\output_filter[3][1] [5]));
   AOI221_X1 i_9_36_51 (.A(n_9_36_46), .B1(n_25), .B2(\buffer[0][3][1] [5]), 
      .C1(\buffer[12][3][1] [5]), .C2(n_27), .ZN(n_9_36_45));
   NAND4_X1 i_9_36_52 (.A1(n_9_36_52), .A2(n_9_36_50), .A3(n_9_36_48), .A4(
      n_9_36_47), .ZN(n_9_36_46));
   AOI22_X1 i_9_36_53 (.A1(\buffer[15][3][1] [5]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][1] [5]), .ZN(n_9_36_47));
   AOI22_X1 i_9_36_54 (.A1(\buffer[10][3][1] [5]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][1] [5]), .ZN(n_9_36_48));
   AOI22_X1 i_9_36_55 (.A1(\buffer[6][3][1] [5]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][1] [5]), .ZN(n_9_36_49));
   AOI22_X1 i_9_36_56 (.A1(\buffer[9][3][1] [5]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][3][1] [5]), .ZN(n_9_36_50));
   AOI22_X1 i_9_36_57 (.A1(\buffer[14][3][1] [5]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][1] [5]), .ZN(n_9_36_51));
   AOI22_X1 i_9_36_58 (.A1(\buffer[11][3][1] [5]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][1] [5]), .ZN(n_9_36_52));
   AOI22_X1 i_9_36_59 (.A1(\buffer[13][3][1] [5]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][1] [5]), .ZN(n_9_36_53));
   NAND4_X1 i_9_36_60 (.A1(n_9_36_62), .A2(n_9_36_60), .A3(n_9_36_58), .A4(
      n_9_36_54), .ZN(\output_filter[3][1] [6]));
   AOI221_X1 i_9_36_61 (.A(n_9_36_55), .B1(n_25), .B2(\buffer[0][3][1] [6]), 
      .C1(\buffer[12][3][1] [6]), .C2(n_27), .ZN(n_9_36_54));
   NAND4_X1 i_9_36_62 (.A1(n_9_36_61), .A2(n_9_36_59), .A3(n_9_36_57), .A4(
      n_9_36_56), .ZN(n_9_36_55));
   AOI22_X1 i_9_36_63 (.A1(\buffer[15][3][1] [6]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][1] [6]), .ZN(n_9_36_56));
   AOI22_X1 i_9_36_64 (.A1(\buffer[10][3][1] [6]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][1] [6]), .ZN(n_9_36_57));
   AOI22_X1 i_9_36_65 (.A1(\buffer[6][3][1] [6]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][1] [6]), .ZN(n_9_36_58));
   AOI22_X1 i_9_36_66 (.A1(\buffer[9][3][1] [6]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][3][1] [6]), .ZN(n_9_36_59));
   AOI22_X1 i_9_36_67 (.A1(\buffer[14][3][1] [6]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][1] [6]), .ZN(n_9_36_60));
   AOI22_X1 i_9_36_68 (.A1(\buffer[11][3][1] [6]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][1] [6]), .ZN(n_9_36_61));
   AOI22_X1 i_9_36_69 (.A1(\buffer[13][3][1] [6]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][1] [6]), .ZN(n_9_36_62));
   NAND4_X1 i_9_36_70 (.A1(n_9_36_71), .A2(n_9_36_69), .A3(n_9_36_67), .A4(
      n_9_36_63), .ZN(\output_filter[3][1] [7]));
   AOI221_X1 i_9_36_71 (.A(n_9_36_64), .B1(n_25), .B2(\buffer[0][3][1] [7]), 
      .C1(\buffer[12][3][1] [7]), .C2(n_27), .ZN(n_9_36_63));
   NAND4_X1 i_9_36_72 (.A1(n_9_36_70), .A2(n_9_36_68), .A3(n_9_36_66), .A4(
      n_9_36_65), .ZN(n_9_36_64));
   AOI22_X1 i_9_36_73 (.A1(\buffer[15][3][1] [7]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][1] [7]), .ZN(n_9_36_65));
   AOI22_X1 i_9_36_74 (.A1(\buffer[10][3][1] [7]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][1] [7]), .ZN(n_9_36_66));
   AOI22_X1 i_9_36_75 (.A1(\buffer[6][3][1] [7]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][1] [7]), .ZN(n_9_36_67));
   AOI22_X1 i_9_36_76 (.A1(\buffer[9][3][1] [7]), .A2(n_20), .B1(n_24), .B2(
      \buffer[2][3][1] [7]), .ZN(n_9_36_68));
   AOI22_X1 i_9_36_77 (.A1(\buffer[14][3][1] [7]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][1] [7]), .ZN(n_9_36_69));
   AOI22_X1 i_9_36_78 (.A1(\buffer[11][3][1] [7]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][1] [7]), .ZN(n_9_36_70));
   AOI22_X1 i_9_36_79 (.A1(\buffer[13][3][1] [7]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][3][1] [7]), .ZN(n_9_36_71));
   NAND4_X1 i_9_36_80 (.A1(n_9_36_80), .A2(n_9_36_78), .A3(n_9_36_76), .A4(
      n_9_36_72), .ZN(\output_filter[3][1] [8]));
   AOI221_X1 i_9_36_81 (.A(n_9_36_73), .B1(n_25), .B2(\buffer[0][3][1] [8]), 
      .C1(\buffer[12][3][1] [8]), .C2(n_27), .ZN(n_9_36_72));
   NAND4_X1 i_9_36_82 (.A1(n_9_36_79), .A2(n_9_36_77), .A3(n_9_36_75), .A4(
      n_9_36_74), .ZN(n_9_36_73));
   AOI22_X1 i_9_36_83 (.A1(\buffer[15][3][1] [8]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][1] [8]), .ZN(n_9_36_74));
   AOI22_X1 i_9_36_84 (.A1(\buffer[10][3][1] [8]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][1] [8]), .ZN(n_9_36_75));
   AOI22_X1 i_9_36_85 (.A1(\buffer[6][3][1] [8]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][1] [8]), .ZN(n_9_36_76));
   AOI22_X1 i_9_36_86 (.A1(\buffer[9][3][1] [8]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][3][1] [8]), .ZN(n_9_36_77));
   AOI22_X1 i_9_36_87 (.A1(\buffer[14][3][1] [8]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][1] [8]), .ZN(n_9_36_78));
   AOI22_X1 i_9_36_88 (.A1(\buffer[11][3][1] [8]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][1] [8]), .ZN(n_9_36_79));
   AOI22_X1 i_9_36_89 (.A1(\buffer[13][3][1] [8]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][1] [8]), .ZN(n_9_36_80));
   NAND4_X1 i_9_36_90 (.A1(n_9_36_89), .A2(n_9_36_87), .A3(n_9_36_85), .A4(
      n_9_36_81), .ZN(\output_filter[3][1] [9]));
   AOI221_X1 i_9_36_91 (.A(n_9_36_82), .B1(n_25), .B2(\buffer[0][3][1] [9]), 
      .C1(\buffer[12][3][1] [9]), .C2(n_27), .ZN(n_9_36_81));
   NAND4_X1 i_9_36_92 (.A1(n_9_36_88), .A2(n_9_36_86), .A3(n_9_36_84), .A4(
      n_9_36_83), .ZN(n_9_36_82));
   AOI22_X1 i_9_36_93 (.A1(\buffer[15][3][1] [9]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][1] [9]), .ZN(n_9_36_83));
   AOI22_X1 i_9_36_94 (.A1(\buffer[10][3][1] [9]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][1] [9]), .ZN(n_9_36_84));
   AOI22_X1 i_9_36_95 (.A1(\buffer[6][3][1] [9]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][1] [9]), .ZN(n_9_36_85));
   AOI22_X1 i_9_36_96 (.A1(\buffer[9][3][1] [9]), .A2(n_20), .B1(n_24), .B2(
      \buffer[2][3][1] [9]), .ZN(n_9_36_86));
   AOI22_X1 i_9_36_97 (.A1(\buffer[14][3][1] [9]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][1] [9]), .ZN(n_9_36_87));
   AOI22_X1 i_9_36_98 (.A1(\buffer[11][3][1] [9]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][1] [9]), .ZN(n_9_36_88));
   AOI22_X1 i_9_36_99 (.A1(\buffer[13][3][1] [9]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][3][1] [9]), .ZN(n_9_36_89));
   NAND4_X1 i_9_36_100 (.A1(n_9_36_98), .A2(n_9_36_96), .A3(n_9_36_94), .A4(
      n_9_36_90), .ZN(\output_filter[3][1] [10]));
   AOI221_X1 i_9_36_101 (.A(n_9_36_91), .B1(n_25), .B2(\buffer[0][3][1] [10]), 
      .C1(\buffer[12][3][1] [10]), .C2(n_27), .ZN(n_9_36_90));
   NAND4_X1 i_9_36_102 (.A1(n_9_36_97), .A2(n_9_36_95), .A3(n_9_36_93), .A4(
      n_9_36_92), .ZN(n_9_36_91));
   AOI22_X1 i_9_36_103 (.A1(\buffer[15][3][1] [10]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][1] [10]), .ZN(n_9_36_92));
   AOI22_X1 i_9_36_104 (.A1(\buffer[10][3][1] [10]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][1] [10]), .ZN(n_9_36_93));
   AOI22_X1 i_9_36_105 (.A1(\buffer[6][3][1] [10]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][1] [10]), .ZN(n_9_36_94));
   AOI22_X1 i_9_36_106 (.A1(\buffer[9][3][1] [10]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][3][1] [10]), .ZN(n_9_36_95));
   AOI22_X1 i_9_36_107 (.A1(\buffer[14][3][1] [10]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][1] [10]), .ZN(n_9_36_96));
   AOI22_X1 i_9_36_108 (.A1(\buffer[11][3][1] [10]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][1] [10]), .ZN(n_9_36_97));
   AOI22_X1 i_9_36_109 (.A1(\buffer[13][3][1] [10]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][1] [10]), .ZN(n_9_36_98));
   NAND4_X1 i_9_36_110 (.A1(n_9_36_107), .A2(n_9_36_105), .A3(n_9_36_103), 
      .A4(n_9_36_99), .ZN(\output_filter[3][1] [11]));
   AOI221_X1 i_9_36_111 (.A(n_9_36_100), .B1(n_25), .B2(\buffer[0][3][1] [11]), 
      .C1(\buffer[12][3][1] [11]), .C2(n_27), .ZN(n_9_36_99));
   NAND4_X1 i_9_36_112 (.A1(n_9_36_106), .A2(n_9_36_104), .A3(n_9_36_102), 
      .A4(n_9_36_101), .ZN(n_9_36_100));
   AOI22_X1 i_9_36_113 (.A1(\buffer[15][3][1] [11]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][1] [11]), .ZN(n_9_36_101));
   AOI22_X1 i_9_36_114 (.A1(\buffer[10][3][1] [11]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][1] [11]), .ZN(n_9_36_102));
   AOI22_X1 i_9_36_115 (.A1(\buffer[6][3][1] [11]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][1] [11]), .ZN(n_9_36_103));
   AOI22_X1 i_9_36_116 (.A1(\buffer[9][3][1] [11]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][3][1] [11]), .ZN(n_9_36_104));
   AOI22_X1 i_9_36_117 (.A1(\buffer[14][3][1] [11]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][1] [11]), .ZN(n_9_36_105));
   AOI22_X1 i_9_36_118 (.A1(\buffer[11][3][1] [11]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][1] [11]), .ZN(n_9_36_106));
   AOI22_X1 i_9_36_119 (.A1(\buffer[13][3][1] [11]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][3][1] [11]), .ZN(n_9_36_107));
   NAND4_X1 i_9_36_120 (.A1(n_9_36_116), .A2(n_9_36_114), .A3(n_9_36_112), 
      .A4(n_9_36_108), .ZN(\output_filter[3][1] [12]));
   AOI221_X1 i_9_36_121 (.A(n_9_36_109), .B1(n_25), .B2(\buffer[0][3][1] [12]), 
      .C1(\buffer[12][3][1] [12]), .C2(n_27), .ZN(n_9_36_108));
   NAND4_X1 i_9_36_122 (.A1(n_9_36_115), .A2(n_9_36_113), .A3(n_9_36_111), 
      .A4(n_9_36_110), .ZN(n_9_36_109));
   AOI22_X1 i_9_36_123 (.A1(\buffer[15][3][1] [12]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][1] [12]), .ZN(n_9_36_110));
   AOI22_X1 i_9_36_124 (.A1(\buffer[10][3][1] [12]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][1] [12]), .ZN(n_9_36_111));
   AOI22_X1 i_9_36_125 (.A1(\buffer[6][3][1] [12]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][1] [12]), .ZN(n_9_36_112));
   AOI22_X1 i_9_36_126 (.A1(\buffer[9][3][1] [12]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][3][1] [12]), .ZN(n_9_36_113));
   AOI22_X1 i_9_36_127 (.A1(\buffer[14][3][1] [12]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][1] [12]), .ZN(n_9_36_114));
   AOI22_X1 i_9_36_128 (.A1(\buffer[11][3][1] [12]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][1] [12]), .ZN(n_9_36_115));
   AOI22_X1 i_9_36_129 (.A1(\buffer[13][3][1] [12]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][1] [12]), .ZN(n_9_36_116));
   NAND4_X1 i_9_36_130 (.A1(n_9_36_125), .A2(n_9_36_123), .A3(n_9_36_121), 
      .A4(n_9_36_117), .ZN(\output_filter[3][1] [13]));
   AOI221_X1 i_9_36_131 (.A(n_9_36_118), .B1(n_25), .B2(\buffer[0][3][1] [13]), 
      .C1(\buffer[12][3][1] [13]), .C2(n_27), .ZN(n_9_36_117));
   NAND4_X1 i_9_36_132 (.A1(n_9_36_124), .A2(n_9_36_122), .A3(n_9_36_120), 
      .A4(n_9_36_119), .ZN(n_9_36_118));
   AOI22_X1 i_9_36_133 (.A1(\buffer[15][3][1] [13]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][1] [13]), .ZN(n_9_36_119));
   AOI22_X1 i_9_36_134 (.A1(\buffer[10][3][1] [13]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][1] [13]), .ZN(n_9_36_120));
   AOI22_X1 i_9_36_135 (.A1(\buffer[6][3][1] [13]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][1] [13]), .ZN(n_9_36_121));
   AOI22_X1 i_9_36_136 (.A1(\buffer[9][3][1] [13]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][3][1] [13]), .ZN(n_9_36_122));
   AOI22_X1 i_9_36_137 (.A1(\buffer[14][3][1] [13]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][1] [13]), .ZN(n_9_36_123));
   AOI22_X1 i_9_36_138 (.A1(\buffer[11][3][1] [13]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][1] [13]), .ZN(n_9_36_124));
   AOI22_X1 i_9_36_139 (.A1(\buffer[13][3][1] [13]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][3][1] [13]), .ZN(n_9_36_125));
   NAND4_X1 i_9_36_140 (.A1(n_9_36_134), .A2(n_9_36_132), .A3(n_9_36_130), 
      .A4(n_9_36_126), .ZN(\output_filter[3][1] [14]));
   AOI221_X1 i_9_36_141 (.A(n_9_36_127), .B1(n_25), .B2(\buffer[0][3][1] [14]), 
      .C1(\buffer[12][3][1] [14]), .C2(n_27), .ZN(n_9_36_126));
   NAND4_X1 i_9_36_142 (.A1(n_9_36_133), .A2(n_9_36_131), .A3(n_9_36_129), 
      .A4(n_9_36_128), .ZN(n_9_36_127));
   AOI22_X1 i_9_36_143 (.A1(\buffer[15][3][1] [14]), .A2(n_22), .B1(n_16), 
      .B2(\buffer[8][3][1] [14]), .ZN(n_9_36_128));
   AOI22_X1 i_9_36_144 (.A1(\buffer[10][3][1] [14]), .A2(n_21), .B1(n_29), 
      .B2(\buffer[7][3][1] [14]), .ZN(n_9_36_129));
   AOI22_X1 i_9_36_145 (.A1(\buffer[6][3][1] [14]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][1] [14]), .ZN(n_9_36_130));
   AOI22_X1 i_9_36_146 (.A1(\buffer[9][3][1] [14]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][3][1] [14]), .ZN(n_9_36_131));
   AOI22_X1 i_9_36_147 (.A1(\buffer[14][3][1] [14]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][1] [14]), .ZN(n_9_36_132));
   AOI22_X1 i_9_36_148 (.A1(\buffer[11][3][1] [14]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][1] [14]), .ZN(n_9_36_133));
   AOI22_X1 i_9_36_149 (.A1(\buffer[13][3][1] [14]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][1] [14]), .ZN(n_9_36_134));
   NAND2_X1 i_9_36_150 (.A1(n_9_36_137), .A2(n_9_36_135), .ZN(
      \output_filter[3][1] [15]));
   AOI221_X1 i_9_36_151 (.A(n_9_36_136), .B1(n_31), .B2(\buffer[3][3][1] [15]), 
      .C1(\buffer[14][3][1] [15]), .C2(n_19), .ZN(n_9_36_135));
   NAND3_X1 i_9_36_152 (.A1(n_9_36_143), .A2(n_9_36_141), .A3(n_9_36_139), 
      .ZN(n_9_36_136));
   AOI221_X1 i_9_36_153 (.A(n_9_36_138), .B1(n_16), .B2(\buffer[8][3][1] [15]), 
      .C1(\buffer[13][3][1] [15]), .C2(n_26), .ZN(n_9_36_137));
   NAND3_X1 i_9_36_154 (.A1(n_9_36_144), .A2(n_9_36_142), .A3(n_9_36_140), 
      .ZN(n_9_36_138));
   AOI22_X1 i_9_36_155 (.A1(\buffer[11][3][1] [15]), .A2(n_17), .B1(n_24), 
      .B2(\buffer[2][3][1] [15]), .ZN(n_9_36_139));
   AOI22_X1 i_9_36_156 (.A1(\buffer[10][3][1] [15]), .A2(n_21), .B1(n_23), 
      .B2(\buffer[1][3][1] [15]), .ZN(n_9_36_140));
   AOI22_X1 i_9_36_157 (.A1(\buffer[6][3][1] [15]), .A2(n_28), .B1(n_18), 
      .B2(\buffer[5][3][1] [15]), .ZN(n_9_36_141));
   AOI22_X1 i_9_36_158 (.A1(\buffer[9][3][1] [15]), .A2(n_20), .B1(n_30), 
      .B2(\buffer[4][3][1] [15]), .ZN(n_9_36_142));
   AOI22_X1 i_9_36_159 (.A1(\buffer[7][3][1] [15]), .A2(n_29), .B1(n_25), 
      .B2(\buffer[0][3][1] [15]), .ZN(n_9_36_143));
   AOI22_X1 i_9_36_160 (.A1(\buffer[15][3][1] [15]), .A2(n_22), .B1(n_27), 
      .B2(\buffer[12][3][1] [15]), .ZN(n_9_36_144));
   NAND4_X1 i_10_35_0 (.A1(n_10_35_8), .A2(n_10_35_6), .A3(n_10_35_4), .A4(
      n_10_35_0), .ZN(\output_filter[3][0] [0]));
   AOI221_X1 i_10_35_1 (.A(n_10_35_1), .B1(n_25), .B2(\buffer[0][3][0] [0]), 
      .C1(\buffer[12][3][0] [0]), .C2(n_27), .ZN(n_10_35_0));
   NAND4_X1 i_10_35_2 (.A1(n_10_35_7), .A2(n_10_35_5), .A3(n_10_35_3), .A4(
      n_10_35_2), .ZN(n_10_35_1));
   AOI22_X1 i_10_35_3 (.A1(\buffer[15][3][0] [0]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][0] [0]), .ZN(n_10_35_2));
   AOI22_X1 i_10_35_4 (.A1(\buffer[10][3][0] [0]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][0] [0]), .ZN(n_10_35_3));
   AOI22_X1 i_10_35_5 (.A1(\buffer[6][3][0] [0]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][0] [0]), .ZN(n_10_35_4));
   AOI22_X1 i_10_35_6 (.A1(\buffer[9][3][0] [0]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][3][0] [0]), .ZN(n_10_35_5));
   AOI22_X1 i_10_35_7 (.A1(\buffer[14][3][0] [0]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][0] [0]), .ZN(n_10_35_6));
   AOI22_X1 i_10_35_8 (.A1(\buffer[11][3][0] [0]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][0] [0]), .ZN(n_10_35_7));
   AOI22_X1 i_10_35_9 (.A1(\buffer[13][3][0] [0]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][0] [0]), .ZN(n_10_35_8));
   NAND4_X1 i_10_35_10 (.A1(n_10_35_17), .A2(n_10_35_15), .A3(n_10_35_13), 
      .A4(n_10_35_9), .ZN(\output_filter[3][0] [1]));
   AOI221_X1 i_10_35_11 (.A(n_10_35_10), .B1(n_25), .B2(\buffer[0][3][0] [1]), 
      .C1(\buffer[12][3][0] [1]), .C2(n_27), .ZN(n_10_35_9));
   NAND4_X1 i_10_35_12 (.A1(n_10_35_16), .A2(n_10_35_14), .A3(n_10_35_12), 
      .A4(n_10_35_11), .ZN(n_10_35_10));
   AOI22_X1 i_10_35_13 (.A1(\buffer[15][3][0] [1]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][0] [1]), .ZN(n_10_35_11));
   AOI22_X1 i_10_35_14 (.A1(\buffer[10][3][0] [1]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][0] [1]), .ZN(n_10_35_12));
   AOI22_X1 i_10_35_15 (.A1(\buffer[6][3][0] [1]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][0] [1]), .ZN(n_10_35_13));
   AOI22_X1 i_10_35_16 (.A1(\buffer[9][3][0] [1]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][3][0] [1]), .ZN(n_10_35_14));
   AOI22_X1 i_10_35_17 (.A1(\buffer[14][3][0] [1]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][0] [1]), .ZN(n_10_35_15));
   AOI22_X1 i_10_35_18 (.A1(\buffer[11][3][0] [1]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][0] [1]), .ZN(n_10_35_16));
   AOI22_X1 i_10_35_19 (.A1(\buffer[13][3][0] [1]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][0] [1]), .ZN(n_10_35_17));
   NAND4_X1 i_10_35_20 (.A1(n_10_35_26), .A2(n_10_35_24), .A3(n_10_35_22), 
      .A4(n_10_35_18), .ZN(\output_filter[3][0] [2]));
   AOI221_X1 i_10_35_21 (.A(n_10_35_19), .B1(n_25), .B2(\buffer[0][3][0] [2]), 
      .C1(\buffer[12][3][0] [2]), .C2(n_27), .ZN(n_10_35_18));
   NAND4_X1 i_10_35_22 (.A1(n_10_35_25), .A2(n_10_35_23), .A3(n_10_35_21), 
      .A4(n_10_35_20), .ZN(n_10_35_19));
   AOI22_X1 i_10_35_23 (.A1(\buffer[15][3][0] [2]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][0] [2]), .ZN(n_10_35_20));
   AOI22_X1 i_10_35_24 (.A1(\buffer[10][3][0] [2]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][0] [2]), .ZN(n_10_35_21));
   AOI22_X1 i_10_35_25 (.A1(\buffer[6][3][0] [2]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][0] [2]), .ZN(n_10_35_22));
   AOI22_X1 i_10_35_26 (.A1(\buffer[9][3][0] [2]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][3][0] [2]), .ZN(n_10_35_23));
   AOI22_X1 i_10_35_27 (.A1(\buffer[14][3][0] [2]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][0] [2]), .ZN(n_10_35_24));
   AOI22_X1 i_10_35_28 (.A1(\buffer[11][3][0] [2]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][0] [2]), .ZN(n_10_35_25));
   AOI22_X1 i_10_35_29 (.A1(\buffer[13][3][0] [2]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][0] [2]), .ZN(n_10_35_26));
   NAND4_X1 i_10_35_30 (.A1(n_10_35_35), .A2(n_10_35_33), .A3(n_10_35_31), 
      .A4(n_10_35_27), .ZN(\output_filter[3][0] [3]));
   AOI221_X1 i_10_35_31 (.A(n_10_35_28), .B1(n_25), .B2(\buffer[0][3][0] [3]), 
      .C1(\buffer[12][3][0] [3]), .C2(n_27), .ZN(n_10_35_27));
   NAND4_X1 i_10_35_32 (.A1(n_10_35_34), .A2(n_10_35_32), .A3(n_10_35_30), 
      .A4(n_10_35_29), .ZN(n_10_35_28));
   AOI22_X1 i_10_35_33 (.A1(\buffer[15][3][0] [3]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][0] [3]), .ZN(n_10_35_29));
   AOI22_X1 i_10_35_34 (.A1(\buffer[10][3][0] [3]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][0] [3]), .ZN(n_10_35_30));
   AOI22_X1 i_10_35_35 (.A1(\buffer[6][3][0] [3]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][0] [3]), .ZN(n_10_35_31));
   AOI22_X1 i_10_35_36 (.A1(\buffer[9][3][0] [3]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][3][0] [3]), .ZN(n_10_35_32));
   AOI22_X1 i_10_35_37 (.A1(\buffer[14][3][0] [3]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][0] [3]), .ZN(n_10_35_33));
   AOI22_X1 i_10_35_38 (.A1(\buffer[11][3][0] [3]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][0] [3]), .ZN(n_10_35_34));
   AOI22_X1 i_10_35_39 (.A1(\buffer[13][3][0] [3]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][0] [3]), .ZN(n_10_35_35));
   NAND4_X1 i_10_35_40 (.A1(n_10_35_44), .A2(n_10_35_42), .A3(n_10_35_40), 
      .A4(n_10_35_36), .ZN(\output_filter[3][0] [4]));
   AOI221_X1 i_10_35_41 (.A(n_10_35_37), .B1(n_25), .B2(\buffer[0][3][0] [4]), 
      .C1(\buffer[12][3][0] [4]), .C2(n_27), .ZN(n_10_35_36));
   NAND4_X1 i_10_35_42 (.A1(n_10_35_43), .A2(n_10_35_41), .A3(n_10_35_39), 
      .A4(n_10_35_38), .ZN(n_10_35_37));
   AOI22_X1 i_10_35_43 (.A1(\buffer[15][3][0] [4]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][0] [4]), .ZN(n_10_35_38));
   AOI22_X1 i_10_35_44 (.A1(\buffer[10][3][0] [4]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][0] [4]), .ZN(n_10_35_39));
   AOI22_X1 i_10_35_45 (.A1(\buffer[6][3][0] [4]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][0] [4]), .ZN(n_10_35_40));
   AOI22_X1 i_10_35_46 (.A1(\buffer[9][3][0] [4]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][3][0] [4]), .ZN(n_10_35_41));
   AOI22_X1 i_10_35_47 (.A1(\buffer[14][3][0] [4]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][0] [4]), .ZN(n_10_35_42));
   AOI22_X1 i_10_35_48 (.A1(\buffer[11][3][0] [4]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][0] [4]), .ZN(n_10_35_43));
   AOI22_X1 i_10_35_49 (.A1(\buffer[13][3][0] [4]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][3][0] [4]), .ZN(n_10_35_44));
   NAND4_X1 i_10_35_50 (.A1(n_10_35_53), .A2(n_10_35_51), .A3(n_10_35_49), 
      .A4(n_10_35_45), .ZN(\output_filter[3][0] [5]));
   AOI221_X1 i_10_35_51 (.A(n_10_35_46), .B1(n_25), .B2(\buffer[0][3][0] [5]), 
      .C1(\buffer[12][3][0] [5]), .C2(n_27), .ZN(n_10_35_45));
   NAND4_X1 i_10_35_52 (.A1(n_10_35_52), .A2(n_10_35_50), .A3(n_10_35_48), 
      .A4(n_10_35_47), .ZN(n_10_35_46));
   AOI22_X1 i_10_35_53 (.A1(\buffer[15][3][0] [5]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][0] [5]), .ZN(n_10_35_47));
   AOI22_X1 i_10_35_54 (.A1(\buffer[10][3][0] [5]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][0] [5]), .ZN(n_10_35_48));
   AOI22_X1 i_10_35_55 (.A1(\buffer[6][3][0] [5]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][0] [5]), .ZN(n_10_35_49));
   AOI22_X1 i_10_35_56 (.A1(\buffer[9][3][0] [5]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][3][0] [5]), .ZN(n_10_35_50));
   AOI22_X1 i_10_35_57 (.A1(\buffer[14][3][0] [5]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][0] [5]), .ZN(n_10_35_51));
   AOI22_X1 i_10_35_58 (.A1(\buffer[11][3][0] [5]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][0] [5]), .ZN(n_10_35_52));
   AOI22_X1 i_10_35_59 (.A1(\buffer[13][3][0] [5]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][0] [5]), .ZN(n_10_35_53));
   NAND4_X1 i_10_35_60 (.A1(n_10_35_62), .A2(n_10_35_60), .A3(n_10_35_58), 
      .A4(n_10_35_54), .ZN(\output_filter[3][0] [6]));
   AOI221_X1 i_10_35_61 (.A(n_10_35_55), .B1(n_25), .B2(\buffer[0][3][0] [6]), 
      .C1(\buffer[12][3][0] [6]), .C2(n_27), .ZN(n_10_35_54));
   NAND4_X1 i_10_35_62 (.A1(n_10_35_61), .A2(n_10_35_59), .A3(n_10_35_57), 
      .A4(n_10_35_56), .ZN(n_10_35_55));
   AOI22_X1 i_10_35_63 (.A1(\buffer[15][3][0] [6]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][0] [6]), .ZN(n_10_35_56));
   AOI22_X1 i_10_35_64 (.A1(\buffer[10][3][0] [6]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][0] [6]), .ZN(n_10_35_57));
   AOI22_X1 i_10_35_65 (.A1(\buffer[6][3][0] [6]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][0] [6]), .ZN(n_10_35_58));
   AOI22_X1 i_10_35_66 (.A1(\buffer[9][3][0] [6]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][3][0] [6]), .ZN(n_10_35_59));
   AOI22_X1 i_10_35_67 (.A1(\buffer[14][3][0] [6]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][0] [6]), .ZN(n_10_35_60));
   AOI22_X1 i_10_35_68 (.A1(\buffer[11][3][0] [6]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][0] [6]), .ZN(n_10_35_61));
   AOI22_X1 i_10_35_69 (.A1(\buffer[13][3][0] [6]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][0] [6]), .ZN(n_10_35_62));
   NAND4_X1 i_10_35_70 (.A1(n_10_35_71), .A2(n_10_35_69), .A3(n_10_35_67), 
      .A4(n_10_35_63), .ZN(\output_filter[3][0] [7]));
   AOI221_X1 i_10_35_71 (.A(n_10_35_64), .B1(n_25), .B2(\buffer[0][3][0] [7]), 
      .C1(\buffer[12][3][0] [7]), .C2(n_27), .ZN(n_10_35_63));
   NAND4_X1 i_10_35_72 (.A1(n_10_35_70), .A2(n_10_35_68), .A3(n_10_35_66), 
      .A4(n_10_35_65), .ZN(n_10_35_64));
   AOI22_X1 i_10_35_73 (.A1(\buffer[15][3][0] [7]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][0] [7]), .ZN(n_10_35_65));
   AOI22_X1 i_10_35_74 (.A1(\buffer[10][3][0] [7]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][0] [7]), .ZN(n_10_35_66));
   AOI22_X1 i_10_35_75 (.A1(\buffer[6][3][0] [7]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][0] [7]), .ZN(n_10_35_67));
   AOI22_X1 i_10_35_76 (.A1(\buffer[9][3][0] [7]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][3][0] [7]), .ZN(n_10_35_68));
   AOI22_X1 i_10_35_77 (.A1(\buffer[14][3][0] [7]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][0] [7]), .ZN(n_10_35_69));
   AOI22_X1 i_10_35_78 (.A1(\buffer[11][3][0] [7]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][0] [7]), .ZN(n_10_35_70));
   AOI22_X1 i_10_35_79 (.A1(\buffer[13][3][0] [7]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][3][0] [7]), .ZN(n_10_35_71));
   NAND4_X1 i_10_35_80 (.A1(n_10_35_80), .A2(n_10_35_78), .A3(n_10_35_76), 
      .A4(n_10_35_72), .ZN(\output_filter[3][0] [8]));
   AOI221_X1 i_10_35_81 (.A(n_10_35_73), .B1(n_25), .B2(\buffer[0][3][0] [8]), 
      .C1(\buffer[12][3][0] [8]), .C2(n_27), .ZN(n_10_35_72));
   NAND4_X1 i_10_35_82 (.A1(n_10_35_79), .A2(n_10_35_77), .A3(n_10_35_75), 
      .A4(n_10_35_74), .ZN(n_10_35_73));
   AOI22_X1 i_10_35_83 (.A1(\buffer[15][3][0] [8]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][0] [8]), .ZN(n_10_35_74));
   AOI22_X1 i_10_35_84 (.A1(\buffer[10][3][0] [8]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][0] [8]), .ZN(n_10_35_75));
   AOI22_X1 i_10_35_85 (.A1(\buffer[6][3][0] [8]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][0] [8]), .ZN(n_10_35_76));
   AOI22_X1 i_10_35_86 (.A1(\buffer[9][3][0] [8]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][3][0] [8]), .ZN(n_10_35_77));
   AOI22_X1 i_10_35_87 (.A1(\buffer[14][3][0] [8]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][0] [8]), .ZN(n_10_35_78));
   AOI22_X1 i_10_35_88 (.A1(\buffer[11][3][0] [8]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][0] [8]), .ZN(n_10_35_79));
   AOI22_X1 i_10_35_89 (.A1(\buffer[13][3][0] [8]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][0] [8]), .ZN(n_10_35_80));
   NAND4_X1 i_10_35_90 (.A1(n_10_35_89), .A2(n_10_35_87), .A3(n_10_35_85), 
      .A4(n_10_35_81), .ZN(\output_filter[3][0] [9]));
   AOI221_X1 i_10_35_91 (.A(n_10_35_82), .B1(n_25), .B2(\buffer[0][3][0] [9]), 
      .C1(\buffer[12][3][0] [9]), .C2(n_27), .ZN(n_10_35_81));
   NAND4_X1 i_10_35_92 (.A1(n_10_35_88), .A2(n_10_35_86), .A3(n_10_35_84), 
      .A4(n_10_35_83), .ZN(n_10_35_82));
   AOI22_X1 i_10_35_93 (.A1(\buffer[15][3][0] [9]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][0] [9]), .ZN(n_10_35_83));
   AOI22_X1 i_10_35_94 (.A1(\buffer[10][3][0] [9]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][0] [9]), .ZN(n_10_35_84));
   AOI22_X1 i_10_35_95 (.A1(\buffer[6][3][0] [9]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][0] [9]), .ZN(n_10_35_85));
   AOI22_X1 i_10_35_96 (.A1(\buffer[9][3][0] [9]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][3][0] [9]), .ZN(n_10_35_86));
   AOI22_X1 i_10_35_97 (.A1(\buffer[14][3][0] [9]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][0] [9]), .ZN(n_10_35_87));
   AOI22_X1 i_10_35_98 (.A1(\buffer[11][3][0] [9]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][0] [9]), .ZN(n_10_35_88));
   AOI22_X1 i_10_35_99 (.A1(\buffer[13][3][0] [9]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][3][0] [9]), .ZN(n_10_35_89));
   NAND4_X1 i_10_35_100 (.A1(n_10_35_98), .A2(n_10_35_96), .A3(n_10_35_94), 
      .A4(n_10_35_90), .ZN(\output_filter[3][0] [10]));
   AOI221_X1 i_10_35_101 (.A(n_10_35_91), .B1(n_25), .B2(\buffer[0][3][0] [10]), 
      .C1(\buffer[12][3][0] [10]), .C2(n_27), .ZN(n_10_35_90));
   NAND4_X1 i_10_35_102 (.A1(n_10_35_97), .A2(n_10_35_95), .A3(n_10_35_93), 
      .A4(n_10_35_92), .ZN(n_10_35_91));
   AOI22_X1 i_10_35_103 (.A1(\buffer[15][3][0] [10]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][0] [10]), .ZN(n_10_35_92));
   AOI22_X1 i_10_35_104 (.A1(\buffer[10][3][0] [10]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][0] [10]), .ZN(n_10_35_93));
   AOI22_X1 i_10_35_105 (.A1(\buffer[6][3][0] [10]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][0] [10]), .ZN(n_10_35_94));
   AOI22_X1 i_10_35_106 (.A1(\buffer[9][3][0] [10]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][3][0] [10]), .ZN(n_10_35_95));
   AOI22_X1 i_10_35_107 (.A1(\buffer[14][3][0] [10]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][0] [10]), .ZN(n_10_35_96));
   AOI22_X1 i_10_35_108 (.A1(\buffer[11][3][0] [10]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][0] [10]), .ZN(n_10_35_97));
   AOI22_X1 i_10_35_109 (.A1(\buffer[13][3][0] [10]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][0] [10]), .ZN(n_10_35_98));
   NAND4_X1 i_10_35_110 (.A1(n_10_35_107), .A2(n_10_35_105), .A3(n_10_35_103), 
      .A4(n_10_35_99), .ZN(\output_filter[3][0] [11]));
   AOI221_X1 i_10_35_111 (.A(n_10_35_100), .B1(n_25), .B2(\buffer[0][3][0] [11]), 
      .C1(\buffer[12][3][0] [11]), .C2(n_27), .ZN(n_10_35_99));
   NAND4_X1 i_10_35_112 (.A1(n_10_35_106), .A2(n_10_35_104), .A3(n_10_35_102), 
      .A4(n_10_35_101), .ZN(n_10_35_100));
   AOI22_X1 i_10_35_113 (.A1(\buffer[15][3][0] [11]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][0] [11]), .ZN(n_10_35_101));
   AOI22_X1 i_10_35_114 (.A1(\buffer[10][3][0] [11]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][0] [11]), .ZN(n_10_35_102));
   AOI22_X1 i_10_35_115 (.A1(\buffer[6][3][0] [11]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][0] [11]), .ZN(n_10_35_103));
   AOI22_X1 i_10_35_116 (.A1(\buffer[9][3][0] [11]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][3][0] [11]), .ZN(n_10_35_104));
   AOI22_X1 i_10_35_117 (.A1(\buffer[14][3][0] [11]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][0] [11]), .ZN(n_10_35_105));
   AOI22_X1 i_10_35_118 (.A1(\buffer[11][3][0] [11]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][0] [11]), .ZN(n_10_35_106));
   AOI22_X1 i_10_35_119 (.A1(\buffer[13][3][0] [11]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][3][0] [11]), .ZN(n_10_35_107));
   NAND4_X1 i_10_35_120 (.A1(n_10_35_116), .A2(n_10_35_114), .A3(n_10_35_112), 
      .A4(n_10_35_108), .ZN(\output_filter[3][0] [12]));
   AOI221_X1 i_10_35_121 (.A(n_10_35_109), .B1(n_25), .B2(\buffer[0][3][0] [12]), 
      .C1(\buffer[12][3][0] [12]), .C2(n_27), .ZN(n_10_35_108));
   NAND4_X1 i_10_35_122 (.A1(n_10_35_115), .A2(n_10_35_113), .A3(n_10_35_111), 
      .A4(n_10_35_110), .ZN(n_10_35_109));
   AOI22_X1 i_10_35_123 (.A1(\buffer[15][3][0] [12]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][0] [12]), .ZN(n_10_35_110));
   AOI22_X1 i_10_35_124 (.A1(\buffer[10][3][0] [12]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][0] [12]), .ZN(n_10_35_111));
   AOI22_X1 i_10_35_125 (.A1(\buffer[6][3][0] [12]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][0] [12]), .ZN(n_10_35_112));
   AOI22_X1 i_10_35_126 (.A1(\buffer[9][3][0] [12]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][3][0] [12]), .ZN(n_10_35_113));
   AOI22_X1 i_10_35_127 (.A1(\buffer[14][3][0] [12]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][0] [12]), .ZN(n_10_35_114));
   AOI22_X1 i_10_35_128 (.A1(\buffer[11][3][0] [12]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][0] [12]), .ZN(n_10_35_115));
   AOI22_X1 i_10_35_129 (.A1(\buffer[13][3][0] [12]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][0] [12]), .ZN(n_10_35_116));
   NAND4_X1 i_10_35_130 (.A1(n_10_35_125), .A2(n_10_35_123), .A3(n_10_35_121), 
      .A4(n_10_35_117), .ZN(\output_filter[3][0] [13]));
   AOI221_X1 i_10_35_131 (.A(n_10_35_118), .B1(n_25), .B2(\buffer[0][3][0] [13]), 
      .C1(\buffer[12][3][0] [13]), .C2(n_27), .ZN(n_10_35_117));
   NAND4_X1 i_10_35_132 (.A1(n_10_35_124), .A2(n_10_35_122), .A3(n_10_35_120), 
      .A4(n_10_35_119), .ZN(n_10_35_118));
   AOI22_X1 i_10_35_133 (.A1(\buffer[15][3][0] [13]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][0] [13]), .ZN(n_10_35_119));
   AOI22_X1 i_10_35_134 (.A1(\buffer[10][3][0] [13]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][0] [13]), .ZN(n_10_35_120));
   AOI22_X1 i_10_35_135 (.A1(\buffer[6][3][0] [13]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][0] [13]), .ZN(n_10_35_121));
   AOI22_X1 i_10_35_136 (.A1(\buffer[9][3][0] [13]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][3][0] [13]), .ZN(n_10_35_122));
   AOI22_X1 i_10_35_137 (.A1(\buffer[14][3][0] [13]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][0] [13]), .ZN(n_10_35_123));
   AOI22_X1 i_10_35_138 (.A1(\buffer[11][3][0] [13]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][0] [13]), .ZN(n_10_35_124));
   AOI22_X1 i_10_35_139 (.A1(\buffer[13][3][0] [13]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][3][0] [13]), .ZN(n_10_35_125));
   NAND4_X1 i_10_35_140 (.A1(n_10_35_134), .A2(n_10_35_132), .A3(n_10_35_130), 
      .A4(n_10_35_126), .ZN(\output_filter[3][0] [14]));
   AOI221_X1 i_10_35_141 (.A(n_10_35_127), .B1(n_25), .B2(\buffer[0][3][0] [14]), 
      .C1(\buffer[12][3][0] [14]), .C2(n_27), .ZN(n_10_35_126));
   NAND4_X1 i_10_35_142 (.A1(n_10_35_133), .A2(n_10_35_131), .A3(n_10_35_129), 
      .A4(n_10_35_128), .ZN(n_10_35_127));
   AOI22_X1 i_10_35_143 (.A1(\buffer[15][3][0] [14]), .A2(n_22), .B1(n_16), 
      .B2(\buffer[8][3][0] [14]), .ZN(n_10_35_128));
   AOI22_X1 i_10_35_144 (.A1(\buffer[10][3][0] [14]), .A2(n_21), .B1(n_29), 
      .B2(\buffer[7][3][0] [14]), .ZN(n_10_35_129));
   AOI22_X1 i_10_35_145 (.A1(\buffer[6][3][0] [14]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][0] [14]), .ZN(n_10_35_130));
   AOI22_X1 i_10_35_146 (.A1(\buffer[9][3][0] [14]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][3][0] [14]), .ZN(n_10_35_131));
   AOI22_X1 i_10_35_147 (.A1(\buffer[14][3][0] [14]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][0] [14]), .ZN(n_10_35_132));
   AOI22_X1 i_10_35_148 (.A1(\buffer[11][3][0] [14]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][0] [14]), .ZN(n_10_35_133));
   AOI22_X1 i_10_35_149 (.A1(\buffer[13][3][0] [14]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][0] [14]), .ZN(n_10_35_134));
   NAND2_X1 i_10_35_150 (.A1(n_10_35_137), .A2(n_10_35_135), .ZN(
      \output_filter[3][0] [15]));
   AOI221_X1 i_10_35_151 (.A(n_10_35_136), .B1(n_31), .B2(\buffer[3][3][0] [15]), 
      .C1(\buffer[14][3][0] [15]), .C2(n_19), .ZN(n_10_35_135));
   NAND3_X1 i_10_35_152 (.A1(n_10_35_143), .A2(n_10_35_141), .A3(n_10_35_139), 
      .ZN(n_10_35_136));
   AOI221_X1 i_10_35_153 (.A(n_10_35_138), .B1(n_16), .B2(\buffer[8][3][0] [15]), 
      .C1(\buffer[13][3][0] [15]), .C2(n_26), .ZN(n_10_35_137));
   NAND3_X1 i_10_35_154 (.A1(n_10_35_144), .A2(n_10_35_142), .A3(n_10_35_140), 
      .ZN(n_10_35_138));
   AOI22_X1 i_10_35_155 (.A1(\buffer[11][3][0] [15]), .A2(n_17), .B1(n_24), 
      .B2(\buffer[2][3][0] [15]), .ZN(n_10_35_139));
   AOI22_X1 i_10_35_156 (.A1(\buffer[10][3][0] [15]), .A2(n_21), .B1(n_23), 
      .B2(\buffer[1][3][0] [15]), .ZN(n_10_35_140));
   AOI22_X1 i_10_35_157 (.A1(\buffer[6][3][0] [15]), .A2(n_28), .B1(n_18), 
      .B2(\buffer[5][3][0] [15]), .ZN(n_10_35_141));
   AOI22_X1 i_10_35_158 (.A1(\buffer[9][3][0] [15]), .A2(n_20), .B1(n_30), 
      .B2(\buffer[4][3][0] [15]), .ZN(n_10_35_142));
   AOI22_X1 i_10_35_159 (.A1(\buffer[7][3][0] [15]), .A2(n_29), .B1(n_25), 
      .B2(\buffer[0][3][0] [15]), .ZN(n_10_35_143));
   AOI22_X1 i_10_35_160 (.A1(\buffer[15][3][0] [15]), .A2(n_22), .B1(n_27), 
      .B2(\buffer[12][3][0] [15]), .ZN(n_10_35_144));
   NAND4_X1 i_11_33_0 (.A1(n_11_33_8), .A2(n_11_33_6), .A3(n_11_33_4), .A4(
      n_11_33_0), .ZN(\output_filter[2][3] [0]));
   AOI221_X1 i_11_33_1 (.A(n_11_33_1), .B1(n_25), .B2(\buffer[0][2][3] [0]), 
      .C1(\buffer[12][2][3] [0]), .C2(n_27), .ZN(n_11_33_0));
   NAND4_X1 i_11_33_2 (.A1(n_11_33_7), .A2(n_11_33_5), .A3(n_11_33_3), .A4(
      n_11_33_2), .ZN(n_11_33_1));
   AOI22_X1 i_11_33_3 (.A1(\buffer[15][2][3] [0]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][3] [0]), .ZN(n_11_33_2));
   AOI22_X1 i_11_33_4 (.A1(\buffer[10][2][3] [0]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][3] [0]), .ZN(n_11_33_3));
   AOI22_X1 i_11_33_5 (.A1(\buffer[6][2][3] [0]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][2][3] [0]), .ZN(n_11_33_4));
   AOI22_X1 i_11_33_6 (.A1(\buffer[9][2][3] [0]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][2][3] [0]), .ZN(n_11_33_5));
   AOI22_X1 i_11_33_7 (.A1(\buffer[14][2][3] [0]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][3] [0]), .ZN(n_11_33_6));
   AOI22_X1 i_11_33_8 (.A1(\buffer[11][2][3] [0]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][3] [0]), .ZN(n_11_33_7));
   AOI22_X1 i_11_33_9 (.A1(\buffer[13][2][3] [0]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][3] [0]), .ZN(n_11_33_8));
   NAND4_X1 i_11_33_10 (.A1(n_11_33_17), .A2(n_11_33_15), .A3(n_11_33_13), 
      .A4(n_11_33_9), .ZN(\output_filter[2][3] [1]));
   AOI221_X1 i_11_33_11 (.A(n_11_33_10), .B1(n_25), .B2(\buffer[0][2][3] [1]), 
      .C1(\buffer[12][2][3] [1]), .C2(n_27), .ZN(n_11_33_9));
   NAND4_X1 i_11_33_12 (.A1(n_11_33_16), .A2(n_11_33_14), .A3(n_11_33_12), 
      .A4(n_11_33_11), .ZN(n_11_33_10));
   AOI22_X1 i_11_33_13 (.A1(\buffer[15][2][3] [1]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][3] [1]), .ZN(n_11_33_11));
   AOI22_X1 i_11_33_14 (.A1(\buffer[10][2][3] [1]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][3] [1]), .ZN(n_11_33_12));
   AOI22_X1 i_11_33_15 (.A1(\buffer[6][2][3] [1]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][3] [1]), .ZN(n_11_33_13));
   AOI22_X1 i_11_33_16 (.A1(\buffer[9][2][3] [1]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][3] [1]), .ZN(n_11_33_14));
   AOI22_X1 i_11_33_17 (.A1(\buffer[14][2][3] [1]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][3] [1]), .ZN(n_11_33_15));
   AOI22_X1 i_11_33_18 (.A1(\buffer[11][2][3] [1]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][3] [1]), .ZN(n_11_33_16));
   AOI22_X1 i_11_33_19 (.A1(\buffer[13][2][3] [1]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][3] [1]), .ZN(n_11_33_17));
   NAND4_X1 i_11_33_20 (.A1(n_11_33_26), .A2(n_11_33_24), .A3(n_11_33_22), 
      .A4(n_11_33_18), .ZN(\output_filter[2][3] [2]));
   AOI221_X1 i_11_33_21 (.A(n_11_33_19), .B1(n_25), .B2(\buffer[0][2][3] [2]), 
      .C1(\buffer[12][2][3] [2]), .C2(n_27), .ZN(n_11_33_18));
   NAND4_X1 i_11_33_22 (.A1(n_11_33_25), .A2(n_11_33_23), .A3(n_11_33_21), 
      .A4(n_11_33_20), .ZN(n_11_33_19));
   AOI22_X1 i_11_33_23 (.A1(\buffer[15][2][3] [2]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][3] [2]), .ZN(n_11_33_20));
   AOI22_X1 i_11_33_24 (.A1(\buffer[10][2][3] [2]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][3] [2]), .ZN(n_11_33_21));
   AOI22_X1 i_11_33_25 (.A1(\buffer[6][2][3] [2]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][3] [2]), .ZN(n_11_33_22));
   AOI22_X1 i_11_33_26 (.A1(\buffer[9][2][3] [2]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][3] [2]), .ZN(n_11_33_23));
   AOI22_X1 i_11_33_27 (.A1(\buffer[14][2][3] [2]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][3] [2]), .ZN(n_11_33_24));
   AOI22_X1 i_11_33_28 (.A1(\buffer[11][2][3] [2]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][3] [2]), .ZN(n_11_33_25));
   AOI22_X1 i_11_33_29 (.A1(\buffer[13][2][3] [2]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][3] [2]), .ZN(n_11_33_26));
   NAND4_X1 i_11_33_30 (.A1(n_11_33_35), .A2(n_11_33_33), .A3(n_11_33_31), 
      .A4(n_11_33_27), .ZN(\output_filter[2][3] [3]));
   AOI221_X1 i_11_33_31 (.A(n_11_33_28), .B1(n_25), .B2(\buffer[0][2][3] [3]), 
      .C1(\buffer[12][2][3] [3]), .C2(n_27), .ZN(n_11_33_27));
   NAND4_X1 i_11_33_32 (.A1(n_11_33_34), .A2(n_11_33_32), .A3(n_11_33_30), 
      .A4(n_11_33_29), .ZN(n_11_33_28));
   AOI22_X1 i_11_33_33 (.A1(\buffer[15][2][3] [3]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][3] [3]), .ZN(n_11_33_29));
   AOI22_X1 i_11_33_34 (.A1(\buffer[10][2][3] [3]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][3] [3]), .ZN(n_11_33_30));
   AOI22_X1 i_11_33_35 (.A1(\buffer[6][2][3] [3]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][3] [3]), .ZN(n_11_33_31));
   AOI22_X1 i_11_33_36 (.A1(\buffer[9][2][3] [3]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][3] [3]), .ZN(n_11_33_32));
   AOI22_X1 i_11_33_37 (.A1(\buffer[14][2][3] [3]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][3] [3]), .ZN(n_11_33_33));
   AOI22_X1 i_11_33_38 (.A1(\buffer[11][2][3] [3]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][3] [3]), .ZN(n_11_33_34));
   AOI22_X1 i_11_33_39 (.A1(\buffer[13][2][3] [3]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][3] [3]), .ZN(n_11_33_35));
   NAND4_X1 i_11_33_40 (.A1(n_11_33_44), .A2(n_11_33_42), .A3(n_11_33_40), 
      .A4(n_11_33_36), .ZN(\output_filter[2][3] [4]));
   AOI221_X1 i_11_33_41 (.A(n_11_33_37), .B1(n_25), .B2(\buffer[0][2][3] [4]), 
      .C1(\buffer[12][2][3] [4]), .C2(n_27), .ZN(n_11_33_36));
   NAND4_X1 i_11_33_42 (.A1(n_11_33_43), .A2(n_11_33_41), .A3(n_11_33_39), 
      .A4(n_11_33_38), .ZN(n_11_33_37));
   AOI22_X1 i_11_33_43 (.A1(\buffer[15][2][3] [4]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][3] [4]), .ZN(n_11_33_38));
   AOI22_X1 i_11_33_44 (.A1(\buffer[10][2][3] [4]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][3] [4]), .ZN(n_11_33_39));
   AOI22_X1 i_11_33_45 (.A1(\buffer[6][2][3] [4]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][3] [4]), .ZN(n_11_33_40));
   AOI22_X1 i_11_33_46 (.A1(\buffer[9][2][3] [4]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][2][3] [4]), .ZN(n_11_33_41));
   AOI22_X1 i_11_33_47 (.A1(\buffer[14][2][3] [4]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][3] [4]), .ZN(n_11_33_42));
   AOI22_X1 i_11_33_48 (.A1(\buffer[11][2][3] [4]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][3] [4]), .ZN(n_11_33_43));
   AOI22_X1 i_11_33_49 (.A1(\buffer[13][2][3] [4]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][2][3] [4]), .ZN(n_11_33_44));
   NAND4_X1 i_11_33_50 (.A1(n_11_33_53), .A2(n_11_33_51), .A3(n_11_33_49), 
      .A4(n_11_33_45), .ZN(\output_filter[2][3] [5]));
   AOI221_X1 i_11_33_51 (.A(n_11_33_46), .B1(n_25), .B2(\buffer[0][2][3] [5]), 
      .C1(\buffer[12][2][3] [5]), .C2(n_27), .ZN(n_11_33_45));
   NAND4_X1 i_11_33_52 (.A1(n_11_33_52), .A2(n_11_33_50), .A3(n_11_33_48), 
      .A4(n_11_33_47), .ZN(n_11_33_46));
   AOI22_X1 i_11_33_53 (.A1(\buffer[15][2][3] [5]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][3] [5]), .ZN(n_11_33_47));
   AOI22_X1 i_11_33_54 (.A1(\buffer[10][2][3] [5]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][3] [5]), .ZN(n_11_33_48));
   AOI22_X1 i_11_33_55 (.A1(\buffer[6][2][3] [5]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][3] [5]), .ZN(n_11_33_49));
   AOI22_X1 i_11_33_56 (.A1(\buffer[9][2][3] [5]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][3] [5]), .ZN(n_11_33_50));
   AOI22_X1 i_11_33_57 (.A1(\buffer[14][2][3] [5]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][3] [5]), .ZN(n_11_33_51));
   AOI22_X1 i_11_33_58 (.A1(\buffer[11][2][3] [5]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][3] [5]), .ZN(n_11_33_52));
   AOI22_X1 i_11_33_59 (.A1(\buffer[13][2][3] [5]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][3] [5]), .ZN(n_11_33_53));
   NAND4_X1 i_11_33_60 (.A1(n_11_33_62), .A2(n_11_33_60), .A3(n_11_33_58), 
      .A4(n_11_33_54), .ZN(\output_filter[2][3] [6]));
   AOI221_X1 i_11_33_61 (.A(n_11_33_55), .B1(n_25), .B2(\buffer[0][2][3] [6]), 
      .C1(\buffer[12][2][3] [6]), .C2(n_27), .ZN(n_11_33_54));
   NAND4_X1 i_11_33_62 (.A1(n_11_33_61), .A2(n_11_33_59), .A3(n_11_33_57), 
      .A4(n_11_33_56), .ZN(n_11_33_55));
   AOI22_X1 i_11_33_63 (.A1(\buffer[15][2][3] [6]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][3] [6]), .ZN(n_11_33_56));
   AOI22_X1 i_11_33_64 (.A1(\buffer[10][2][3] [6]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][3] [6]), .ZN(n_11_33_57));
   AOI22_X1 i_11_33_65 (.A1(\buffer[6][2][3] [6]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][3] [6]), .ZN(n_11_33_58));
   AOI22_X1 i_11_33_66 (.A1(\buffer[9][2][3] [6]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][3] [6]), .ZN(n_11_33_59));
   AOI22_X1 i_11_33_67 (.A1(\buffer[14][2][3] [6]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][3] [6]), .ZN(n_11_33_60));
   AOI22_X1 i_11_33_68 (.A1(\buffer[11][2][3] [6]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][3] [6]), .ZN(n_11_33_61));
   AOI22_X1 i_11_33_69 (.A1(\buffer[13][2][3] [6]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][3] [6]), .ZN(n_11_33_62));
   NAND4_X1 i_11_33_70 (.A1(n_11_33_71), .A2(n_11_33_69), .A3(n_11_33_67), 
      .A4(n_11_33_63), .ZN(\output_filter[2][3] [7]));
   AOI221_X1 i_11_33_71 (.A(n_11_33_64), .B1(n_25), .B2(\buffer[0][2][3] [7]), 
      .C1(\buffer[12][2][3] [7]), .C2(n_27), .ZN(n_11_33_63));
   NAND4_X1 i_11_33_72 (.A1(n_11_33_70), .A2(n_11_33_68), .A3(n_11_33_66), 
      .A4(n_11_33_65), .ZN(n_11_33_64));
   AOI22_X1 i_11_33_73 (.A1(\buffer[15][2][3] [7]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][3] [7]), .ZN(n_11_33_65));
   AOI22_X1 i_11_33_74 (.A1(\buffer[10][2][3] [7]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][3] [7]), .ZN(n_11_33_66));
   AOI22_X1 i_11_33_75 (.A1(\buffer[6][2][3] [7]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][3] [7]), .ZN(n_11_33_67));
   AOI22_X1 i_11_33_76 (.A1(\buffer[9][2][3] [7]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][2][3] [7]), .ZN(n_11_33_68));
   AOI22_X1 i_11_33_77 (.A1(\buffer[14][2][3] [7]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][3] [7]), .ZN(n_11_33_69));
   AOI22_X1 i_11_33_78 (.A1(\buffer[11][2][3] [7]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][3] [7]), .ZN(n_11_33_70));
   AOI22_X1 i_11_33_79 (.A1(\buffer[13][2][3] [7]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][2][3] [7]), .ZN(n_11_33_71));
   NAND4_X1 i_11_33_80 (.A1(n_11_33_80), .A2(n_11_33_78), .A3(n_11_33_76), 
      .A4(n_11_33_72), .ZN(\output_filter[2][3] [8]));
   AOI221_X1 i_11_33_81 (.A(n_11_33_73), .B1(n_25), .B2(\buffer[0][2][3] [8]), 
      .C1(\buffer[12][2][3] [8]), .C2(n_27), .ZN(n_11_33_72));
   NAND4_X1 i_11_33_82 (.A1(n_11_33_79), .A2(n_11_33_77), .A3(n_11_33_75), 
      .A4(n_11_33_74), .ZN(n_11_33_73));
   AOI22_X1 i_11_33_83 (.A1(\buffer[15][2][3] [8]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][3] [8]), .ZN(n_11_33_74));
   AOI22_X1 i_11_33_84 (.A1(\buffer[10][2][3] [8]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][3] [8]), .ZN(n_11_33_75));
   AOI22_X1 i_11_33_85 (.A1(\buffer[6][2][3] [8]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][3] [8]), .ZN(n_11_33_76));
   AOI22_X1 i_11_33_86 (.A1(\buffer[9][2][3] [8]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][3] [8]), .ZN(n_11_33_77));
   AOI22_X1 i_11_33_87 (.A1(\buffer[14][2][3] [8]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][3] [8]), .ZN(n_11_33_78));
   AOI22_X1 i_11_33_88 (.A1(\buffer[11][2][3] [8]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][3] [8]), .ZN(n_11_33_79));
   AOI22_X1 i_11_33_89 (.A1(\buffer[13][2][3] [8]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][3] [8]), .ZN(n_11_33_80));
   NAND4_X1 i_11_33_90 (.A1(n_11_33_89), .A2(n_11_33_87), .A3(n_11_33_85), 
      .A4(n_11_33_81), .ZN(\output_filter[2][3] [9]));
   AOI221_X1 i_11_33_91 (.A(n_11_33_82), .B1(n_25), .B2(\buffer[0][2][3] [9]), 
      .C1(\buffer[12][2][3] [9]), .C2(n_27), .ZN(n_11_33_81));
   NAND4_X1 i_11_33_92 (.A1(n_11_33_88), .A2(n_11_33_86), .A3(n_11_33_84), 
      .A4(n_11_33_83), .ZN(n_11_33_82));
   AOI22_X1 i_11_33_93 (.A1(\buffer[15][2][3] [9]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][3] [9]), .ZN(n_11_33_83));
   AOI22_X1 i_11_33_94 (.A1(\buffer[10][2][3] [9]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][3] [9]), .ZN(n_11_33_84));
   AOI22_X1 i_11_33_95 (.A1(\buffer[6][2][3] [9]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][3] [9]), .ZN(n_11_33_85));
   AOI22_X1 i_11_33_96 (.A1(\buffer[9][2][3] [9]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][2][3] [9]), .ZN(n_11_33_86));
   AOI22_X1 i_11_33_97 (.A1(\buffer[14][2][3] [9]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][3] [9]), .ZN(n_11_33_87));
   AOI22_X1 i_11_33_98 (.A1(\buffer[11][2][3] [9]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][3] [9]), .ZN(n_11_33_88));
   AOI22_X1 i_11_33_99 (.A1(\buffer[13][2][3] [9]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][2][3] [9]), .ZN(n_11_33_89));
   NAND4_X1 i_11_33_100 (.A1(n_11_33_98), .A2(n_11_33_96), .A3(n_11_33_94), 
      .A4(n_11_33_90), .ZN(\output_filter[2][3] [10]));
   AOI221_X1 i_11_33_101 (.A(n_11_33_91), .B1(n_25), .B2(\buffer[0][2][3] [10]), 
      .C1(\buffer[12][2][3] [10]), .C2(n_27), .ZN(n_11_33_90));
   NAND4_X1 i_11_33_102 (.A1(n_11_33_97), .A2(n_11_33_95), .A3(n_11_33_93), 
      .A4(n_11_33_92), .ZN(n_11_33_91));
   AOI22_X1 i_11_33_103 (.A1(\buffer[15][2][3] [10]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][3] [10]), .ZN(n_11_33_92));
   AOI22_X1 i_11_33_104 (.A1(\buffer[10][2][3] [10]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][3] [10]), .ZN(n_11_33_93));
   AOI22_X1 i_11_33_105 (.A1(\buffer[6][2][3] [10]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][3] [10]), .ZN(n_11_33_94));
   AOI22_X1 i_11_33_106 (.A1(\buffer[9][2][3] [10]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][3] [10]), .ZN(n_11_33_95));
   AOI22_X1 i_11_33_107 (.A1(\buffer[14][2][3] [10]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][3] [10]), .ZN(n_11_33_96));
   AOI22_X1 i_11_33_108 (.A1(\buffer[11][2][3] [10]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][3] [10]), .ZN(n_11_33_97));
   AOI22_X1 i_11_33_109 (.A1(\buffer[13][2][3] [10]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][3] [10]), .ZN(n_11_33_98));
   NAND4_X1 i_11_33_110 (.A1(n_11_33_107), .A2(n_11_33_105), .A3(n_11_33_103), 
      .A4(n_11_33_99), .ZN(\output_filter[2][3] [11]));
   AOI221_X1 i_11_33_111 (.A(n_11_33_100), .B1(n_25), .B2(\buffer[0][2][3] [11]), 
      .C1(\buffer[12][2][3] [11]), .C2(n_27), .ZN(n_11_33_99));
   NAND4_X1 i_11_33_112 (.A1(n_11_33_106), .A2(n_11_33_104), .A3(n_11_33_102), 
      .A4(n_11_33_101), .ZN(n_11_33_100));
   AOI22_X1 i_11_33_113 (.A1(\buffer[15][2][3] [11]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][3] [11]), .ZN(n_11_33_101));
   AOI22_X1 i_11_33_114 (.A1(\buffer[10][2][3] [11]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][3] [11]), .ZN(n_11_33_102));
   AOI22_X1 i_11_33_115 (.A1(\buffer[6][2][3] [11]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][3] [11]), .ZN(n_11_33_103));
   AOI22_X1 i_11_33_116 (.A1(\buffer[9][2][3] [11]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][2][3] [11]), .ZN(n_11_33_104));
   AOI22_X1 i_11_33_117 (.A1(\buffer[14][2][3] [11]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][3] [11]), .ZN(n_11_33_105));
   AOI22_X1 i_11_33_118 (.A1(\buffer[11][2][3] [11]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][3] [11]), .ZN(n_11_33_106));
   AOI22_X1 i_11_33_119 (.A1(\buffer[13][2][3] [11]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][2][3] [11]), .ZN(n_11_33_107));
   NAND4_X1 i_11_33_120 (.A1(n_11_33_116), .A2(n_11_33_114), .A3(n_11_33_112), 
      .A4(n_11_33_108), .ZN(\output_filter[2][3] [12]));
   AOI221_X1 i_11_33_121 (.A(n_11_33_109), .B1(n_25), .B2(\buffer[0][2][3] [12]), 
      .C1(\buffer[12][2][3] [12]), .C2(n_27), .ZN(n_11_33_108));
   NAND4_X1 i_11_33_122 (.A1(n_11_33_115), .A2(n_11_33_113), .A3(n_11_33_111), 
      .A4(n_11_33_110), .ZN(n_11_33_109));
   AOI22_X1 i_11_33_123 (.A1(\buffer[15][2][3] [12]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][3] [12]), .ZN(n_11_33_110));
   AOI22_X1 i_11_33_124 (.A1(\buffer[10][2][3] [12]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][3] [12]), .ZN(n_11_33_111));
   AOI22_X1 i_11_33_125 (.A1(\buffer[6][2][3] [12]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][3] [12]), .ZN(n_11_33_112));
   AOI22_X1 i_11_33_126 (.A1(\buffer[9][2][3] [12]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][3] [12]), .ZN(n_11_33_113));
   AOI22_X1 i_11_33_127 (.A1(\buffer[14][2][3] [12]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][3] [12]), .ZN(n_11_33_114));
   AOI22_X1 i_11_33_128 (.A1(\buffer[11][2][3] [12]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][3] [12]), .ZN(n_11_33_115));
   AOI22_X1 i_11_33_129 (.A1(\buffer[13][2][3] [12]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][3] [12]), .ZN(n_11_33_116));
   NAND4_X1 i_11_33_130 (.A1(n_11_33_125), .A2(n_11_33_123), .A3(n_11_33_121), 
      .A4(n_11_33_117), .ZN(\output_filter[2][3] [13]));
   AOI221_X1 i_11_33_131 (.A(n_11_33_118), .B1(n_25), .B2(\buffer[0][2][3] [13]), 
      .C1(\buffer[12][2][3] [13]), .C2(n_27), .ZN(n_11_33_117));
   NAND4_X1 i_11_33_132 (.A1(n_11_33_124), .A2(n_11_33_122), .A3(n_11_33_120), 
      .A4(n_11_33_119), .ZN(n_11_33_118));
   AOI22_X1 i_11_33_133 (.A1(\buffer[15][2][3] [13]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][3] [13]), .ZN(n_11_33_119));
   AOI22_X1 i_11_33_134 (.A1(\buffer[10][2][3] [13]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][3] [13]), .ZN(n_11_33_120));
   AOI22_X1 i_11_33_135 (.A1(\buffer[6][2][3] [13]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][3] [13]), .ZN(n_11_33_121));
   AOI22_X1 i_11_33_136 (.A1(\buffer[9][2][3] [13]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][2][3] [13]), .ZN(n_11_33_122));
   AOI22_X1 i_11_33_137 (.A1(\buffer[14][2][3] [13]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][3] [13]), .ZN(n_11_33_123));
   AOI22_X1 i_11_33_138 (.A1(\buffer[11][2][3] [13]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][3] [13]), .ZN(n_11_33_124));
   AOI22_X1 i_11_33_139 (.A1(\buffer[13][2][3] [13]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][2][3] [13]), .ZN(n_11_33_125));
   NAND4_X1 i_11_33_140 (.A1(n_11_33_134), .A2(n_11_33_132), .A3(n_11_33_130), 
      .A4(n_11_33_126), .ZN(\output_filter[2][3] [14]));
   AOI221_X1 i_11_33_141 (.A(n_11_33_127), .B1(n_25), .B2(\buffer[0][2][3] [14]), 
      .C1(\buffer[12][2][3] [14]), .C2(n_27), .ZN(n_11_33_126));
   NAND4_X1 i_11_33_142 (.A1(n_11_33_133), .A2(n_11_33_131), .A3(n_11_33_129), 
      .A4(n_11_33_128), .ZN(n_11_33_127));
   AOI22_X1 i_11_33_143 (.A1(\buffer[15][2][3] [14]), .A2(n_22), .B1(n_16), 
      .B2(\buffer[8][2][3] [14]), .ZN(n_11_33_128));
   AOI22_X1 i_11_33_144 (.A1(\buffer[10][2][3] [14]), .A2(n_21), .B1(n_29), 
      .B2(\buffer[7][2][3] [14]), .ZN(n_11_33_129));
   AOI22_X1 i_11_33_145 (.A1(\buffer[6][2][3] [14]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][3] [14]), .ZN(n_11_33_130));
   AOI22_X1 i_11_33_146 (.A1(\buffer[9][2][3] [14]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][3] [14]), .ZN(n_11_33_131));
   AOI22_X1 i_11_33_147 (.A1(\buffer[14][2][3] [14]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][3] [14]), .ZN(n_11_33_132));
   AOI22_X1 i_11_33_148 (.A1(\buffer[11][2][3] [14]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][3] [14]), .ZN(n_11_33_133));
   AOI22_X1 i_11_33_149 (.A1(\buffer[13][2][3] [14]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][3] [14]), .ZN(n_11_33_134));
   NAND2_X1 i_11_33_150 (.A1(n_11_33_137), .A2(n_11_33_135), .ZN(
      \output_filter[2][3] [15]));
   AOI221_X1 i_11_33_151 (.A(n_11_33_136), .B1(n_31), .B2(\buffer[3][2][3] [15]), 
      .C1(\buffer[14][2][3] [15]), .C2(n_19), .ZN(n_11_33_135));
   NAND3_X1 i_11_33_152 (.A1(n_11_33_143), .A2(n_11_33_141), .A3(n_11_33_139), 
      .ZN(n_11_33_136));
   AOI221_X1 i_11_33_153 (.A(n_11_33_138), .B1(n_16), .B2(\buffer[8][2][3] [15]), 
      .C1(\buffer[13][2][3] [15]), .C2(n_26), .ZN(n_11_33_137));
   NAND3_X1 i_11_33_154 (.A1(n_11_33_144), .A2(n_11_33_142), .A3(n_11_33_140), 
      .ZN(n_11_33_138));
   AOI22_X1 i_11_33_155 (.A1(\buffer[11][2][3] [15]), .A2(n_17), .B1(n_24), 
      .B2(\buffer[2][2][3] [15]), .ZN(n_11_33_139));
   AOI22_X1 i_11_33_156 (.A1(\buffer[10][2][3] [15]), .A2(n_21), .B1(n_23), 
      .B2(\buffer[1][2][3] [15]), .ZN(n_11_33_140));
   AOI22_X1 i_11_33_157 (.A1(\buffer[6][2][3] [15]), .A2(n_28), .B1(n_18), 
      .B2(\buffer[5][2][3] [15]), .ZN(n_11_33_141));
   AOI22_X1 i_11_33_158 (.A1(\buffer[9][2][3] [15]), .A2(n_20), .B1(n_30), 
      .B2(\buffer[4][2][3] [15]), .ZN(n_11_33_142));
   AOI22_X1 i_11_33_159 (.A1(\buffer[7][2][3] [15]), .A2(n_29), .B1(n_25), 
      .B2(\buffer[0][2][3] [15]), .ZN(n_11_33_143));
   AOI22_X1 i_11_33_160 (.A1(\buffer[15][2][3] [15]), .A2(n_22), .B1(n_27), 
      .B2(\buffer[12][2][3] [15]), .ZN(n_11_33_144));
   NAND4_X1 i_12_32_0 (.A1(n_12_32_8), .A2(n_12_32_6), .A3(n_12_32_4), .A4(
      n_12_32_0), .ZN(\output_filter[2][2] [0]));
   AOI221_X1 i_12_32_1 (.A(n_12_32_1), .B1(n_25), .B2(\buffer[0][2][2] [0]), 
      .C1(\buffer[12][2][2] [0]), .C2(n_27), .ZN(n_12_32_0));
   NAND4_X1 i_12_32_2 (.A1(n_12_32_7), .A2(n_12_32_5), .A3(n_12_32_3), .A4(
      n_12_32_2), .ZN(n_12_32_1));
   AOI22_X1 i_12_32_3 (.A1(\buffer[15][2][2] [0]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][2] [0]), .ZN(n_12_32_2));
   AOI22_X1 i_12_32_4 (.A1(\buffer[10][2][2] [0]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][2] [0]), .ZN(n_12_32_3));
   AOI22_X1 i_12_32_5 (.A1(\buffer[6][2][2] [0]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][2][2] [0]), .ZN(n_12_32_4));
   AOI22_X1 i_12_32_6 (.A1(\buffer[9][2][2] [0]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][2][2] [0]), .ZN(n_12_32_5));
   AOI22_X1 i_12_32_7 (.A1(\buffer[14][2][2] [0]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][2] [0]), .ZN(n_12_32_6));
   AOI22_X1 i_12_32_8 (.A1(\buffer[11][2][2] [0]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][2] [0]), .ZN(n_12_32_7));
   AOI22_X1 i_12_32_9 (.A1(\buffer[13][2][2] [0]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][2] [0]), .ZN(n_12_32_8));
   NAND4_X1 i_12_32_10 (.A1(n_12_32_17), .A2(n_12_32_15), .A3(n_12_32_13), 
      .A4(n_12_32_9), .ZN(\output_filter[2][2] [1]));
   AOI221_X1 i_12_32_11 (.A(n_12_32_10), .B1(n_25), .B2(\buffer[0][2][2] [1]), 
      .C1(\buffer[12][2][2] [1]), .C2(n_27), .ZN(n_12_32_9));
   NAND4_X1 i_12_32_12 (.A1(n_12_32_16), .A2(n_12_32_14), .A3(n_12_32_12), 
      .A4(n_12_32_11), .ZN(n_12_32_10));
   AOI22_X1 i_12_32_13 (.A1(\buffer[15][2][2] [1]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][2] [1]), .ZN(n_12_32_11));
   AOI22_X1 i_12_32_14 (.A1(\buffer[10][2][2] [1]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][2] [1]), .ZN(n_12_32_12));
   AOI22_X1 i_12_32_15 (.A1(\buffer[6][2][2] [1]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][2] [1]), .ZN(n_12_32_13));
   AOI22_X1 i_12_32_16 (.A1(\buffer[9][2][2] [1]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][2] [1]), .ZN(n_12_32_14));
   AOI22_X1 i_12_32_17 (.A1(\buffer[14][2][2] [1]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][2] [1]), .ZN(n_12_32_15));
   AOI22_X1 i_12_32_18 (.A1(\buffer[11][2][2] [1]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][2] [1]), .ZN(n_12_32_16));
   AOI22_X1 i_12_32_19 (.A1(\buffer[13][2][2] [1]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][2] [1]), .ZN(n_12_32_17));
   NAND4_X1 i_12_32_20 (.A1(n_12_32_26), .A2(n_12_32_24), .A3(n_12_32_22), 
      .A4(n_12_32_18), .ZN(\output_filter[2][2] [2]));
   AOI221_X1 i_12_32_21 (.A(n_12_32_19), .B1(n_25), .B2(\buffer[0][2][2] [2]), 
      .C1(\buffer[12][2][2] [2]), .C2(n_27), .ZN(n_12_32_18));
   NAND4_X1 i_12_32_22 (.A1(n_12_32_25), .A2(n_12_32_23), .A3(n_12_32_21), 
      .A4(n_12_32_20), .ZN(n_12_32_19));
   AOI22_X1 i_12_32_23 (.A1(\buffer[15][2][2] [2]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][2] [2]), .ZN(n_12_32_20));
   AOI22_X1 i_12_32_24 (.A1(\buffer[10][2][2] [2]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][2] [2]), .ZN(n_12_32_21));
   AOI22_X1 i_12_32_25 (.A1(\buffer[6][2][2] [2]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][2] [2]), .ZN(n_12_32_22));
   AOI22_X1 i_12_32_26 (.A1(\buffer[9][2][2] [2]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][2] [2]), .ZN(n_12_32_23));
   AOI22_X1 i_12_32_27 (.A1(\buffer[14][2][2] [2]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][2] [2]), .ZN(n_12_32_24));
   AOI22_X1 i_12_32_28 (.A1(\buffer[11][2][2] [2]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][2] [2]), .ZN(n_12_32_25));
   AOI22_X1 i_12_32_29 (.A1(\buffer[13][2][2] [2]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][2] [2]), .ZN(n_12_32_26));
   NAND4_X1 i_12_32_30 (.A1(n_12_32_35), .A2(n_12_32_33), .A3(n_12_32_31), 
      .A4(n_12_32_27), .ZN(\output_filter[2][2] [3]));
   AOI221_X1 i_12_32_31 (.A(n_12_32_28), .B1(n_25), .B2(\buffer[0][2][2] [3]), 
      .C1(\buffer[12][2][2] [3]), .C2(n_27), .ZN(n_12_32_27));
   NAND4_X1 i_12_32_32 (.A1(n_12_32_34), .A2(n_12_32_32), .A3(n_12_32_30), 
      .A4(n_12_32_29), .ZN(n_12_32_28));
   AOI22_X1 i_12_32_33 (.A1(\buffer[15][2][2] [3]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][2] [3]), .ZN(n_12_32_29));
   AOI22_X1 i_12_32_34 (.A1(\buffer[10][2][2] [3]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][2] [3]), .ZN(n_12_32_30));
   AOI22_X1 i_12_32_35 (.A1(\buffer[6][2][2] [3]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][2] [3]), .ZN(n_12_32_31));
   AOI22_X1 i_12_32_36 (.A1(\buffer[9][2][2] [3]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][2] [3]), .ZN(n_12_32_32));
   AOI22_X1 i_12_32_37 (.A1(\buffer[14][2][2] [3]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][2] [3]), .ZN(n_12_32_33));
   AOI22_X1 i_12_32_38 (.A1(\buffer[11][2][2] [3]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][2] [3]), .ZN(n_12_32_34));
   AOI22_X1 i_12_32_39 (.A1(\buffer[13][2][2] [3]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][2] [3]), .ZN(n_12_32_35));
   NAND4_X1 i_12_32_40 (.A1(n_12_32_44), .A2(n_12_32_42), .A3(n_12_32_40), 
      .A4(n_12_32_36), .ZN(\output_filter[2][2] [4]));
   AOI221_X1 i_12_32_41 (.A(n_12_32_37), .B1(n_25), .B2(\buffer[0][2][2] [4]), 
      .C1(\buffer[12][2][2] [4]), .C2(n_27), .ZN(n_12_32_36));
   NAND4_X1 i_12_32_42 (.A1(n_12_32_43), .A2(n_12_32_41), .A3(n_12_32_39), 
      .A4(n_12_32_38), .ZN(n_12_32_37));
   AOI22_X1 i_12_32_43 (.A1(\buffer[15][2][2] [4]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][2] [4]), .ZN(n_12_32_38));
   AOI22_X1 i_12_32_44 (.A1(\buffer[10][2][2] [4]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][2] [4]), .ZN(n_12_32_39));
   AOI22_X1 i_12_32_45 (.A1(\buffer[6][2][2] [4]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][2] [4]), .ZN(n_12_32_40));
   AOI22_X1 i_12_32_46 (.A1(\buffer[9][2][2] [4]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][2][2] [4]), .ZN(n_12_32_41));
   AOI22_X1 i_12_32_47 (.A1(\buffer[14][2][2] [4]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][2] [4]), .ZN(n_12_32_42));
   AOI22_X1 i_12_32_48 (.A1(\buffer[11][2][2] [4]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][2] [4]), .ZN(n_12_32_43));
   AOI22_X1 i_12_32_49 (.A1(\buffer[13][2][2] [4]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][2][2] [4]), .ZN(n_12_32_44));
   NAND4_X1 i_12_32_50 (.A1(n_12_32_53), .A2(n_12_32_51), .A3(n_12_32_49), 
      .A4(n_12_32_45), .ZN(\output_filter[2][2] [5]));
   AOI221_X1 i_12_32_51 (.A(n_12_32_46), .B1(n_25), .B2(\buffer[0][2][2] [5]), 
      .C1(\buffer[12][2][2] [5]), .C2(n_27), .ZN(n_12_32_45));
   NAND4_X1 i_12_32_52 (.A1(n_12_32_52), .A2(n_12_32_50), .A3(n_12_32_48), 
      .A4(n_12_32_47), .ZN(n_12_32_46));
   AOI22_X1 i_12_32_53 (.A1(\buffer[15][2][2] [5]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][2] [5]), .ZN(n_12_32_47));
   AOI22_X1 i_12_32_54 (.A1(\buffer[10][2][2] [5]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][2] [5]), .ZN(n_12_32_48));
   AOI22_X1 i_12_32_55 (.A1(\buffer[6][2][2] [5]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][2] [5]), .ZN(n_12_32_49));
   AOI22_X1 i_12_32_56 (.A1(\buffer[9][2][2] [5]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][2] [5]), .ZN(n_12_32_50));
   AOI22_X1 i_12_32_57 (.A1(\buffer[14][2][2] [5]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][2] [5]), .ZN(n_12_32_51));
   AOI22_X1 i_12_32_58 (.A1(\buffer[11][2][2] [5]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][2] [5]), .ZN(n_12_32_52));
   AOI22_X1 i_12_32_59 (.A1(\buffer[13][2][2] [5]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][2] [5]), .ZN(n_12_32_53));
   NAND4_X1 i_12_32_60 (.A1(n_12_32_62), .A2(n_12_32_60), .A3(n_12_32_58), 
      .A4(n_12_32_54), .ZN(\output_filter[2][2] [6]));
   AOI221_X1 i_12_32_61 (.A(n_12_32_55), .B1(n_25), .B2(\buffer[0][2][2] [6]), 
      .C1(\buffer[12][2][2] [6]), .C2(n_27), .ZN(n_12_32_54));
   NAND4_X1 i_12_32_62 (.A1(n_12_32_61), .A2(n_12_32_59), .A3(n_12_32_57), 
      .A4(n_12_32_56), .ZN(n_12_32_55));
   AOI22_X1 i_12_32_63 (.A1(\buffer[15][2][2] [6]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][2] [6]), .ZN(n_12_32_56));
   AOI22_X1 i_12_32_64 (.A1(\buffer[10][2][2] [6]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][2] [6]), .ZN(n_12_32_57));
   AOI22_X1 i_12_32_65 (.A1(\buffer[6][2][2] [6]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][2] [6]), .ZN(n_12_32_58));
   AOI22_X1 i_12_32_66 (.A1(\buffer[9][2][2] [6]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][2] [6]), .ZN(n_12_32_59));
   AOI22_X1 i_12_32_67 (.A1(\buffer[14][2][2] [6]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][2] [6]), .ZN(n_12_32_60));
   AOI22_X1 i_12_32_68 (.A1(\buffer[11][2][2] [6]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][2] [6]), .ZN(n_12_32_61));
   AOI22_X1 i_12_32_69 (.A1(\buffer[13][2][2] [6]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][2] [6]), .ZN(n_12_32_62));
   NAND4_X1 i_12_32_70 (.A1(n_12_32_71), .A2(n_12_32_69), .A3(n_12_32_67), 
      .A4(n_12_32_63), .ZN(\output_filter[2][2] [7]));
   AOI221_X1 i_12_32_71 (.A(n_12_32_64), .B1(n_25), .B2(\buffer[0][2][2] [7]), 
      .C1(\buffer[12][2][2] [7]), .C2(n_27), .ZN(n_12_32_63));
   NAND4_X1 i_12_32_72 (.A1(n_12_32_70), .A2(n_12_32_68), .A3(n_12_32_66), 
      .A4(n_12_32_65), .ZN(n_12_32_64));
   AOI22_X1 i_12_32_73 (.A1(\buffer[15][2][2] [7]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][2] [7]), .ZN(n_12_32_65));
   AOI22_X1 i_12_32_74 (.A1(\buffer[10][2][2] [7]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][2] [7]), .ZN(n_12_32_66));
   AOI22_X1 i_12_32_75 (.A1(\buffer[6][2][2] [7]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][2] [7]), .ZN(n_12_32_67));
   AOI22_X1 i_12_32_76 (.A1(\buffer[9][2][2] [7]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][2][2] [7]), .ZN(n_12_32_68));
   AOI22_X1 i_12_32_77 (.A1(\buffer[14][2][2] [7]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][2] [7]), .ZN(n_12_32_69));
   AOI22_X1 i_12_32_78 (.A1(\buffer[11][2][2] [7]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][2] [7]), .ZN(n_12_32_70));
   AOI22_X1 i_12_32_79 (.A1(\buffer[13][2][2] [7]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][2][2] [7]), .ZN(n_12_32_71));
   NAND4_X1 i_12_32_80 (.A1(n_12_32_80), .A2(n_12_32_78), .A3(n_12_32_76), 
      .A4(n_12_32_72), .ZN(\output_filter[2][2] [8]));
   AOI221_X1 i_12_32_81 (.A(n_12_32_73), .B1(n_25), .B2(\buffer[0][2][2] [8]), 
      .C1(\buffer[12][2][2] [8]), .C2(n_27), .ZN(n_12_32_72));
   NAND4_X1 i_12_32_82 (.A1(n_12_32_79), .A2(n_12_32_77), .A3(n_12_32_75), 
      .A4(n_12_32_74), .ZN(n_12_32_73));
   AOI22_X1 i_12_32_83 (.A1(\buffer[15][2][2] [8]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][2] [8]), .ZN(n_12_32_74));
   AOI22_X1 i_12_32_84 (.A1(\buffer[10][2][2] [8]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][2] [8]), .ZN(n_12_32_75));
   AOI22_X1 i_12_32_85 (.A1(\buffer[6][2][2] [8]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][2] [8]), .ZN(n_12_32_76));
   AOI22_X1 i_12_32_86 (.A1(\buffer[9][2][2] [8]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][2] [8]), .ZN(n_12_32_77));
   AOI22_X1 i_12_32_87 (.A1(\buffer[14][2][2] [8]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][2] [8]), .ZN(n_12_32_78));
   AOI22_X1 i_12_32_88 (.A1(\buffer[11][2][2] [8]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][2] [8]), .ZN(n_12_32_79));
   AOI22_X1 i_12_32_89 (.A1(\buffer[13][2][2] [8]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][2] [8]), .ZN(n_12_32_80));
   NAND4_X1 i_12_32_90 (.A1(n_12_32_89), .A2(n_12_32_87), .A3(n_12_32_85), 
      .A4(n_12_32_81), .ZN(\output_filter[2][2] [9]));
   AOI221_X1 i_12_32_91 (.A(n_12_32_82), .B1(n_25), .B2(\buffer[0][2][2] [9]), 
      .C1(\buffer[12][2][2] [9]), .C2(n_27), .ZN(n_12_32_81));
   NAND4_X1 i_12_32_92 (.A1(n_12_32_88), .A2(n_12_32_86), .A3(n_12_32_84), 
      .A4(n_12_32_83), .ZN(n_12_32_82));
   AOI22_X1 i_12_32_93 (.A1(\buffer[15][2][2] [9]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][2] [9]), .ZN(n_12_32_83));
   AOI22_X1 i_12_32_94 (.A1(\buffer[10][2][2] [9]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][2] [9]), .ZN(n_12_32_84));
   AOI22_X1 i_12_32_95 (.A1(\buffer[6][2][2] [9]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][2] [9]), .ZN(n_12_32_85));
   AOI22_X1 i_12_32_96 (.A1(\buffer[9][2][2] [9]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][2][2] [9]), .ZN(n_12_32_86));
   AOI22_X1 i_12_32_97 (.A1(\buffer[14][2][2] [9]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][2] [9]), .ZN(n_12_32_87));
   AOI22_X1 i_12_32_98 (.A1(\buffer[11][2][2] [9]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][2] [9]), .ZN(n_12_32_88));
   AOI22_X1 i_12_32_99 (.A1(\buffer[13][2][2] [9]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][2][2] [9]), .ZN(n_12_32_89));
   NAND4_X1 i_12_32_100 (.A1(n_12_32_98), .A2(n_12_32_96), .A3(n_12_32_94), 
      .A4(n_12_32_90), .ZN(\output_filter[2][2] [10]));
   AOI221_X1 i_12_32_101 (.A(n_12_32_91), .B1(n_25), .B2(\buffer[0][2][2] [10]), 
      .C1(\buffer[12][2][2] [10]), .C2(n_27), .ZN(n_12_32_90));
   NAND4_X1 i_12_32_102 (.A1(n_12_32_97), .A2(n_12_32_95), .A3(n_12_32_93), 
      .A4(n_12_32_92), .ZN(n_12_32_91));
   AOI22_X1 i_12_32_103 (.A1(\buffer[15][2][2] [10]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][2] [10]), .ZN(n_12_32_92));
   AOI22_X1 i_12_32_104 (.A1(\buffer[10][2][2] [10]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][2] [10]), .ZN(n_12_32_93));
   AOI22_X1 i_12_32_105 (.A1(\buffer[6][2][2] [10]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][2] [10]), .ZN(n_12_32_94));
   AOI22_X1 i_12_32_106 (.A1(\buffer[9][2][2] [10]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][2] [10]), .ZN(n_12_32_95));
   AOI22_X1 i_12_32_107 (.A1(\buffer[14][2][2] [10]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][2] [10]), .ZN(n_12_32_96));
   AOI22_X1 i_12_32_108 (.A1(\buffer[11][2][2] [10]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][2] [10]), .ZN(n_12_32_97));
   AOI22_X1 i_12_32_109 (.A1(\buffer[13][2][2] [10]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][2] [10]), .ZN(n_12_32_98));
   NAND4_X1 i_12_32_110 (.A1(n_12_32_107), .A2(n_12_32_105), .A3(n_12_32_103), 
      .A4(n_12_32_99), .ZN(\output_filter[2][2] [11]));
   AOI221_X1 i_12_32_111 (.A(n_12_32_100), .B1(n_25), .B2(\buffer[0][2][2] [11]), 
      .C1(\buffer[12][2][2] [11]), .C2(n_27), .ZN(n_12_32_99));
   NAND4_X1 i_12_32_112 (.A1(n_12_32_106), .A2(n_12_32_104), .A3(n_12_32_102), 
      .A4(n_12_32_101), .ZN(n_12_32_100));
   AOI22_X1 i_12_32_113 (.A1(\buffer[15][2][2] [11]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][2] [11]), .ZN(n_12_32_101));
   AOI22_X1 i_12_32_114 (.A1(\buffer[10][2][2] [11]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][2] [11]), .ZN(n_12_32_102));
   AOI22_X1 i_12_32_115 (.A1(\buffer[6][2][2] [11]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][2] [11]), .ZN(n_12_32_103));
   AOI22_X1 i_12_32_116 (.A1(\buffer[9][2][2] [11]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][2][2] [11]), .ZN(n_12_32_104));
   AOI22_X1 i_12_32_117 (.A1(\buffer[14][2][2] [11]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][2] [11]), .ZN(n_12_32_105));
   AOI22_X1 i_12_32_118 (.A1(\buffer[11][2][2] [11]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][2] [11]), .ZN(n_12_32_106));
   AOI22_X1 i_12_32_119 (.A1(\buffer[13][2][2] [11]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][2][2] [11]), .ZN(n_12_32_107));
   NAND4_X1 i_12_32_120 (.A1(n_12_32_116), .A2(n_12_32_114), .A3(n_12_32_112), 
      .A4(n_12_32_108), .ZN(\output_filter[2][2] [12]));
   AOI221_X1 i_12_32_121 (.A(n_12_32_109), .B1(n_25), .B2(\buffer[0][2][2] [12]), 
      .C1(\buffer[12][2][2] [12]), .C2(n_27), .ZN(n_12_32_108));
   NAND4_X1 i_12_32_122 (.A1(n_12_32_115), .A2(n_12_32_113), .A3(n_12_32_111), 
      .A4(n_12_32_110), .ZN(n_12_32_109));
   AOI22_X1 i_12_32_123 (.A1(\buffer[15][2][2] [12]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][2] [12]), .ZN(n_12_32_110));
   AOI22_X1 i_12_32_124 (.A1(\buffer[10][2][2] [12]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][2] [12]), .ZN(n_12_32_111));
   AOI22_X1 i_12_32_125 (.A1(\buffer[6][2][2] [12]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][2] [12]), .ZN(n_12_32_112));
   AOI22_X1 i_12_32_126 (.A1(\buffer[9][2][2] [12]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][2] [12]), .ZN(n_12_32_113));
   AOI22_X1 i_12_32_127 (.A1(\buffer[14][2][2] [12]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][2] [12]), .ZN(n_12_32_114));
   AOI22_X1 i_12_32_128 (.A1(\buffer[11][2][2] [12]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][2] [12]), .ZN(n_12_32_115));
   AOI22_X1 i_12_32_129 (.A1(\buffer[13][2][2] [12]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][2] [12]), .ZN(n_12_32_116));
   NAND4_X1 i_12_32_130 (.A1(n_12_32_125), .A2(n_12_32_123), .A3(n_12_32_121), 
      .A4(n_12_32_117), .ZN(\output_filter[2][2] [13]));
   AOI221_X1 i_12_32_131 (.A(n_12_32_118), .B1(n_25), .B2(\buffer[0][2][2] [13]), 
      .C1(\buffer[12][2][2] [13]), .C2(n_27), .ZN(n_12_32_117));
   NAND4_X1 i_12_32_132 (.A1(n_12_32_124), .A2(n_12_32_122), .A3(n_12_32_120), 
      .A4(n_12_32_119), .ZN(n_12_32_118));
   AOI22_X1 i_12_32_133 (.A1(\buffer[15][2][2] [13]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][2] [13]), .ZN(n_12_32_119));
   AOI22_X1 i_12_32_134 (.A1(\buffer[10][2][2] [13]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][2] [13]), .ZN(n_12_32_120));
   AOI22_X1 i_12_32_135 (.A1(\buffer[6][2][2] [13]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][2] [13]), .ZN(n_12_32_121));
   AOI22_X1 i_12_32_136 (.A1(\buffer[9][2][2] [13]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][2][2] [13]), .ZN(n_12_32_122));
   AOI22_X1 i_12_32_137 (.A1(\buffer[14][2][2] [13]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][2] [13]), .ZN(n_12_32_123));
   AOI22_X1 i_12_32_138 (.A1(\buffer[11][2][2] [13]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][2] [13]), .ZN(n_12_32_124));
   AOI22_X1 i_12_32_139 (.A1(\buffer[13][2][2] [13]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][2][2] [13]), .ZN(n_12_32_125));
   NAND4_X1 i_12_32_140 (.A1(n_12_32_134), .A2(n_12_32_132), .A3(n_12_32_130), 
      .A4(n_12_32_126), .ZN(\output_filter[2][2] [14]));
   AOI221_X1 i_12_32_141 (.A(n_12_32_127), .B1(n_25), .B2(\buffer[0][2][2] [14]), 
      .C1(\buffer[12][2][2] [14]), .C2(n_27), .ZN(n_12_32_126));
   NAND4_X1 i_12_32_142 (.A1(n_12_32_133), .A2(n_12_32_131), .A3(n_12_32_129), 
      .A4(n_12_32_128), .ZN(n_12_32_127));
   AOI22_X1 i_12_32_143 (.A1(\buffer[15][2][2] [14]), .A2(n_22), .B1(n_16), 
      .B2(\buffer[8][2][2] [14]), .ZN(n_12_32_128));
   AOI22_X1 i_12_32_144 (.A1(\buffer[10][2][2] [14]), .A2(n_21), .B1(n_29), 
      .B2(\buffer[7][2][2] [14]), .ZN(n_12_32_129));
   AOI22_X1 i_12_32_145 (.A1(\buffer[6][2][2] [14]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][2] [14]), .ZN(n_12_32_130));
   AOI22_X1 i_12_32_146 (.A1(\buffer[9][2][2] [14]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][2] [14]), .ZN(n_12_32_131));
   AOI22_X1 i_12_32_147 (.A1(\buffer[14][2][2] [14]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][2] [14]), .ZN(n_12_32_132));
   AOI22_X1 i_12_32_148 (.A1(\buffer[11][2][2] [14]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][2] [14]), .ZN(n_12_32_133));
   AOI22_X1 i_12_32_149 (.A1(\buffer[13][2][2] [14]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][2] [14]), .ZN(n_12_32_134));
   NAND2_X1 i_12_32_150 (.A1(n_12_32_137), .A2(n_12_32_135), .ZN(
      \output_filter[2][2] [15]));
   AOI221_X1 i_12_32_151 (.A(n_12_32_136), .B1(n_31), .B2(\buffer[3][2][2] [15]), 
      .C1(\buffer[14][2][2] [15]), .C2(n_19), .ZN(n_12_32_135));
   NAND3_X1 i_12_32_152 (.A1(n_12_32_143), .A2(n_12_32_141), .A3(n_12_32_139), 
      .ZN(n_12_32_136));
   AOI221_X1 i_12_32_153 (.A(n_12_32_138), .B1(n_16), .B2(\buffer[8][2][2] [15]), 
      .C1(\buffer[13][2][2] [15]), .C2(n_26), .ZN(n_12_32_137));
   NAND3_X1 i_12_32_154 (.A1(n_12_32_144), .A2(n_12_32_142), .A3(n_12_32_140), 
      .ZN(n_12_32_138));
   AOI22_X1 i_12_32_155 (.A1(\buffer[11][2][2] [15]), .A2(n_17), .B1(n_24), 
      .B2(\buffer[2][2][2] [15]), .ZN(n_12_32_139));
   AOI22_X1 i_12_32_156 (.A1(\buffer[10][2][2] [15]), .A2(n_21), .B1(n_23), 
      .B2(\buffer[1][2][2] [15]), .ZN(n_12_32_140));
   AOI22_X1 i_12_32_157 (.A1(\buffer[6][2][2] [15]), .A2(n_28), .B1(n_18), 
      .B2(\buffer[5][2][2] [15]), .ZN(n_12_32_141));
   AOI22_X1 i_12_32_158 (.A1(\buffer[9][2][2] [15]), .A2(n_20), .B1(n_30), 
      .B2(\buffer[4][2][2] [15]), .ZN(n_12_32_142));
   AOI22_X1 i_12_32_159 (.A1(\buffer[7][2][2] [15]), .A2(n_29), .B1(n_25), 
      .B2(\buffer[0][2][2] [15]), .ZN(n_12_32_143));
   AOI22_X1 i_12_32_160 (.A1(\buffer[15][2][2] [15]), .A2(n_22), .B1(n_27), 
      .B2(\buffer[12][2][2] [15]), .ZN(n_12_32_144));
   NAND4_X1 i_13_31_0 (.A1(n_13_31_8), .A2(n_13_31_6), .A3(n_13_31_4), .A4(
      n_13_31_0), .ZN(\output_filter[2][1] [0]));
   AOI221_X1 i_13_31_1 (.A(n_13_31_1), .B1(n_25), .B2(\buffer[0][2][1] [0]), 
      .C1(\buffer[12][2][1] [0]), .C2(n_27), .ZN(n_13_31_0));
   NAND4_X1 i_13_31_2 (.A1(n_13_31_7), .A2(n_13_31_5), .A3(n_13_31_3), .A4(
      n_13_31_2), .ZN(n_13_31_1));
   AOI22_X1 i_13_31_3 (.A1(\buffer[15][2][1] [0]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][1] [0]), .ZN(n_13_31_2));
   AOI22_X1 i_13_31_4 (.A1(\buffer[10][2][1] [0]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][1] [0]), .ZN(n_13_31_3));
   AOI22_X1 i_13_31_5 (.A1(\buffer[6][2][1] [0]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][2][1] [0]), .ZN(n_13_31_4));
   AOI22_X1 i_13_31_6 (.A1(\buffer[9][2][1] [0]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][2][1] [0]), .ZN(n_13_31_5));
   AOI22_X1 i_13_31_7 (.A1(\buffer[14][2][1] [0]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][1] [0]), .ZN(n_13_31_6));
   AOI22_X1 i_13_31_8 (.A1(\buffer[11][2][1] [0]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][1] [0]), .ZN(n_13_31_7));
   AOI22_X1 i_13_31_9 (.A1(\buffer[13][2][1] [0]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][1] [0]), .ZN(n_13_31_8));
   NAND4_X1 i_13_31_10 (.A1(n_13_31_17), .A2(n_13_31_15), .A3(n_13_31_13), 
      .A4(n_13_31_9), .ZN(\output_filter[2][1] [1]));
   AOI221_X1 i_13_31_11 (.A(n_13_31_10), .B1(n_25), .B2(\buffer[0][2][1] [1]), 
      .C1(\buffer[12][2][1] [1]), .C2(n_27), .ZN(n_13_31_9));
   NAND4_X1 i_13_31_12 (.A1(n_13_31_16), .A2(n_13_31_14), .A3(n_13_31_12), 
      .A4(n_13_31_11), .ZN(n_13_31_10));
   AOI22_X1 i_13_31_13 (.A1(\buffer[15][2][1] [1]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][1] [1]), .ZN(n_13_31_11));
   AOI22_X1 i_13_31_14 (.A1(\buffer[10][2][1] [1]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][1] [1]), .ZN(n_13_31_12));
   AOI22_X1 i_13_31_15 (.A1(\buffer[6][2][1] [1]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][1] [1]), .ZN(n_13_31_13));
   AOI22_X1 i_13_31_16 (.A1(\buffer[9][2][1] [1]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][1] [1]), .ZN(n_13_31_14));
   AOI22_X1 i_13_31_17 (.A1(\buffer[14][2][1] [1]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][1] [1]), .ZN(n_13_31_15));
   AOI22_X1 i_13_31_18 (.A1(\buffer[11][2][1] [1]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][1] [1]), .ZN(n_13_31_16));
   AOI22_X1 i_13_31_19 (.A1(\buffer[13][2][1] [1]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][1] [1]), .ZN(n_13_31_17));
   NAND4_X1 i_13_31_20 (.A1(n_13_31_26), .A2(n_13_31_24), .A3(n_13_31_22), 
      .A4(n_13_31_18), .ZN(\output_filter[2][1] [2]));
   AOI221_X1 i_13_31_21 (.A(n_13_31_19), .B1(n_25), .B2(\buffer[0][2][1] [2]), 
      .C1(\buffer[12][2][1] [2]), .C2(n_27), .ZN(n_13_31_18));
   NAND4_X1 i_13_31_22 (.A1(n_13_31_25), .A2(n_13_31_23), .A3(n_13_31_21), 
      .A4(n_13_31_20), .ZN(n_13_31_19));
   AOI22_X1 i_13_31_23 (.A1(\buffer[15][2][1] [2]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][1] [2]), .ZN(n_13_31_20));
   AOI22_X1 i_13_31_24 (.A1(\buffer[10][2][1] [2]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][1] [2]), .ZN(n_13_31_21));
   AOI22_X1 i_13_31_25 (.A1(\buffer[6][2][1] [2]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][1] [2]), .ZN(n_13_31_22));
   AOI22_X1 i_13_31_26 (.A1(\buffer[9][2][1] [2]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][1] [2]), .ZN(n_13_31_23));
   AOI22_X1 i_13_31_27 (.A1(\buffer[14][2][1] [2]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][1] [2]), .ZN(n_13_31_24));
   AOI22_X1 i_13_31_28 (.A1(\buffer[11][2][1] [2]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][1] [2]), .ZN(n_13_31_25));
   AOI22_X1 i_13_31_29 (.A1(\buffer[13][2][1] [2]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][1] [2]), .ZN(n_13_31_26));
   NAND4_X1 i_13_31_30 (.A1(n_13_31_35), .A2(n_13_31_33), .A3(n_13_31_31), 
      .A4(n_13_31_27), .ZN(\output_filter[2][1] [3]));
   AOI221_X1 i_13_31_31 (.A(n_13_31_28), .B1(n_25), .B2(\buffer[0][2][1] [3]), 
      .C1(\buffer[12][2][1] [3]), .C2(n_27), .ZN(n_13_31_27));
   NAND4_X1 i_13_31_32 (.A1(n_13_31_34), .A2(n_13_31_32), .A3(n_13_31_30), 
      .A4(n_13_31_29), .ZN(n_13_31_28));
   AOI22_X1 i_13_31_33 (.A1(\buffer[15][2][1] [3]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][1] [3]), .ZN(n_13_31_29));
   AOI22_X1 i_13_31_34 (.A1(\buffer[10][2][1] [3]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][1] [3]), .ZN(n_13_31_30));
   AOI22_X1 i_13_31_35 (.A1(\buffer[6][2][1] [3]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][1] [3]), .ZN(n_13_31_31));
   AOI22_X1 i_13_31_36 (.A1(\buffer[9][2][1] [3]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][1] [3]), .ZN(n_13_31_32));
   AOI22_X1 i_13_31_37 (.A1(\buffer[14][2][1] [3]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][1] [3]), .ZN(n_13_31_33));
   AOI22_X1 i_13_31_38 (.A1(\buffer[11][2][1] [3]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][1] [3]), .ZN(n_13_31_34));
   AOI22_X1 i_13_31_39 (.A1(\buffer[13][2][1] [3]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][1] [3]), .ZN(n_13_31_35));
   NAND4_X1 i_13_31_40 (.A1(n_13_31_44), .A2(n_13_31_42), .A3(n_13_31_40), 
      .A4(n_13_31_36), .ZN(\output_filter[2][1] [4]));
   AOI221_X1 i_13_31_41 (.A(n_13_31_37), .B1(n_25), .B2(\buffer[0][2][1] [4]), 
      .C1(\buffer[12][2][1] [4]), .C2(n_27), .ZN(n_13_31_36));
   NAND4_X1 i_13_31_42 (.A1(n_13_31_43), .A2(n_13_31_41), .A3(n_13_31_39), 
      .A4(n_13_31_38), .ZN(n_13_31_37));
   AOI22_X1 i_13_31_43 (.A1(\buffer[15][2][1] [4]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][1] [4]), .ZN(n_13_31_38));
   AOI22_X1 i_13_31_44 (.A1(\buffer[10][2][1] [4]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][1] [4]), .ZN(n_13_31_39));
   AOI22_X1 i_13_31_45 (.A1(\buffer[6][2][1] [4]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][1] [4]), .ZN(n_13_31_40));
   AOI22_X1 i_13_31_46 (.A1(\buffer[9][2][1] [4]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][2][1] [4]), .ZN(n_13_31_41));
   AOI22_X1 i_13_31_47 (.A1(\buffer[14][2][1] [4]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][1] [4]), .ZN(n_13_31_42));
   AOI22_X1 i_13_31_48 (.A1(\buffer[11][2][1] [4]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][1] [4]), .ZN(n_13_31_43));
   AOI22_X1 i_13_31_49 (.A1(\buffer[13][2][1] [4]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][2][1] [4]), .ZN(n_13_31_44));
   NAND4_X1 i_13_31_50 (.A1(n_13_31_53), .A2(n_13_31_51), .A3(n_13_31_49), 
      .A4(n_13_31_45), .ZN(\output_filter[2][1] [5]));
   AOI221_X1 i_13_31_51 (.A(n_13_31_46), .B1(n_25), .B2(\buffer[0][2][1] [5]), 
      .C1(\buffer[12][2][1] [5]), .C2(n_27), .ZN(n_13_31_45));
   NAND4_X1 i_13_31_52 (.A1(n_13_31_52), .A2(n_13_31_50), .A3(n_13_31_48), 
      .A4(n_13_31_47), .ZN(n_13_31_46));
   AOI22_X1 i_13_31_53 (.A1(\buffer[15][2][1] [5]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][1] [5]), .ZN(n_13_31_47));
   AOI22_X1 i_13_31_54 (.A1(\buffer[10][2][1] [5]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][1] [5]), .ZN(n_13_31_48));
   AOI22_X1 i_13_31_55 (.A1(\buffer[6][2][1] [5]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][1] [5]), .ZN(n_13_31_49));
   AOI22_X1 i_13_31_56 (.A1(\buffer[9][2][1] [5]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][1] [5]), .ZN(n_13_31_50));
   AOI22_X1 i_13_31_57 (.A1(\buffer[14][2][1] [5]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][1] [5]), .ZN(n_13_31_51));
   AOI22_X1 i_13_31_58 (.A1(\buffer[11][2][1] [5]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][1] [5]), .ZN(n_13_31_52));
   AOI22_X1 i_13_31_59 (.A1(\buffer[13][2][1] [5]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][1] [5]), .ZN(n_13_31_53));
   NAND4_X1 i_13_31_60 (.A1(n_13_31_62), .A2(n_13_31_60), .A3(n_13_31_58), 
      .A4(n_13_31_54), .ZN(\output_filter[2][1] [6]));
   AOI221_X1 i_13_31_61 (.A(n_13_31_55), .B1(n_25), .B2(\buffer[0][2][1] [6]), 
      .C1(\buffer[12][2][1] [6]), .C2(n_27), .ZN(n_13_31_54));
   NAND4_X1 i_13_31_62 (.A1(n_13_31_61), .A2(n_13_31_59), .A3(n_13_31_57), 
      .A4(n_13_31_56), .ZN(n_13_31_55));
   AOI22_X1 i_13_31_63 (.A1(\buffer[15][2][1] [6]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][1] [6]), .ZN(n_13_31_56));
   AOI22_X1 i_13_31_64 (.A1(\buffer[10][2][1] [6]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][1] [6]), .ZN(n_13_31_57));
   AOI22_X1 i_13_31_65 (.A1(\buffer[6][2][1] [6]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][1] [6]), .ZN(n_13_31_58));
   AOI22_X1 i_13_31_66 (.A1(\buffer[9][2][1] [6]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][1] [6]), .ZN(n_13_31_59));
   AOI22_X1 i_13_31_67 (.A1(\buffer[14][2][1] [6]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][1] [6]), .ZN(n_13_31_60));
   AOI22_X1 i_13_31_68 (.A1(\buffer[11][2][1] [6]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][1] [6]), .ZN(n_13_31_61));
   AOI22_X1 i_13_31_69 (.A1(\buffer[13][2][1] [6]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][1] [6]), .ZN(n_13_31_62));
   NAND4_X1 i_13_31_70 (.A1(n_13_31_71), .A2(n_13_31_69), .A3(n_13_31_67), 
      .A4(n_13_31_63), .ZN(\output_filter[2][1] [7]));
   AOI221_X1 i_13_31_71 (.A(n_13_31_64), .B1(n_25), .B2(\buffer[0][2][1] [7]), 
      .C1(\buffer[12][2][1] [7]), .C2(n_27), .ZN(n_13_31_63));
   NAND4_X1 i_13_31_72 (.A1(n_13_31_70), .A2(n_13_31_68), .A3(n_13_31_66), 
      .A4(n_13_31_65), .ZN(n_13_31_64));
   AOI22_X1 i_13_31_73 (.A1(\buffer[15][2][1] [7]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][1] [7]), .ZN(n_13_31_65));
   AOI22_X1 i_13_31_74 (.A1(\buffer[10][2][1] [7]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][1] [7]), .ZN(n_13_31_66));
   AOI22_X1 i_13_31_75 (.A1(\buffer[6][2][1] [7]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][1] [7]), .ZN(n_13_31_67));
   AOI22_X1 i_13_31_76 (.A1(\buffer[9][2][1] [7]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][2][1] [7]), .ZN(n_13_31_68));
   AOI22_X1 i_13_31_77 (.A1(\buffer[14][2][1] [7]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][1] [7]), .ZN(n_13_31_69));
   AOI22_X1 i_13_31_78 (.A1(\buffer[11][2][1] [7]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][1] [7]), .ZN(n_13_31_70));
   AOI22_X1 i_13_31_79 (.A1(\buffer[13][2][1] [7]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][2][1] [7]), .ZN(n_13_31_71));
   NAND4_X1 i_13_31_80 (.A1(n_13_31_80), .A2(n_13_31_78), .A3(n_13_31_76), 
      .A4(n_13_31_72), .ZN(\output_filter[2][1] [8]));
   AOI221_X1 i_13_31_81 (.A(n_13_31_73), .B1(n_25), .B2(\buffer[0][2][1] [8]), 
      .C1(\buffer[12][2][1] [8]), .C2(n_27), .ZN(n_13_31_72));
   NAND4_X1 i_13_31_82 (.A1(n_13_31_79), .A2(n_13_31_77), .A3(n_13_31_75), 
      .A4(n_13_31_74), .ZN(n_13_31_73));
   AOI22_X1 i_13_31_83 (.A1(\buffer[15][2][1] [8]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][1] [8]), .ZN(n_13_31_74));
   AOI22_X1 i_13_31_84 (.A1(\buffer[10][2][1] [8]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][1] [8]), .ZN(n_13_31_75));
   AOI22_X1 i_13_31_85 (.A1(\buffer[6][2][1] [8]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][1] [8]), .ZN(n_13_31_76));
   AOI22_X1 i_13_31_86 (.A1(\buffer[9][2][1] [8]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][1] [8]), .ZN(n_13_31_77));
   AOI22_X1 i_13_31_87 (.A1(\buffer[14][2][1] [8]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][1] [8]), .ZN(n_13_31_78));
   AOI22_X1 i_13_31_88 (.A1(\buffer[11][2][1] [8]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][1] [8]), .ZN(n_13_31_79));
   AOI22_X1 i_13_31_89 (.A1(\buffer[13][2][1] [8]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][1] [8]), .ZN(n_13_31_80));
   NAND4_X1 i_13_31_90 (.A1(n_13_31_89), .A2(n_13_31_87), .A3(n_13_31_85), 
      .A4(n_13_31_81), .ZN(\output_filter[2][1] [9]));
   AOI221_X1 i_13_31_91 (.A(n_13_31_82), .B1(n_25), .B2(\buffer[0][2][1] [9]), 
      .C1(\buffer[12][2][1] [9]), .C2(n_27), .ZN(n_13_31_81));
   NAND4_X1 i_13_31_92 (.A1(n_13_31_88), .A2(n_13_31_86), .A3(n_13_31_84), 
      .A4(n_13_31_83), .ZN(n_13_31_82));
   AOI22_X1 i_13_31_93 (.A1(\buffer[15][2][1] [9]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][1] [9]), .ZN(n_13_31_83));
   AOI22_X1 i_13_31_94 (.A1(\buffer[10][2][1] [9]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][1] [9]), .ZN(n_13_31_84));
   AOI22_X1 i_13_31_95 (.A1(\buffer[6][2][1] [9]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][1] [9]), .ZN(n_13_31_85));
   AOI22_X1 i_13_31_96 (.A1(\buffer[9][2][1] [9]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][2][1] [9]), .ZN(n_13_31_86));
   AOI22_X1 i_13_31_97 (.A1(\buffer[14][2][1] [9]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][1] [9]), .ZN(n_13_31_87));
   AOI22_X1 i_13_31_98 (.A1(\buffer[11][2][1] [9]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][1] [9]), .ZN(n_13_31_88));
   AOI22_X1 i_13_31_99 (.A1(\buffer[13][2][1] [9]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][2][1] [9]), .ZN(n_13_31_89));
   NAND4_X1 i_13_31_100 (.A1(n_13_31_98), .A2(n_13_31_96), .A3(n_13_31_94), 
      .A4(n_13_31_90), .ZN(\output_filter[2][1] [10]));
   AOI221_X1 i_13_31_101 (.A(n_13_31_91), .B1(n_25), .B2(\buffer[0][2][1] [10]), 
      .C1(\buffer[12][2][1] [10]), .C2(n_27), .ZN(n_13_31_90));
   NAND4_X1 i_13_31_102 (.A1(n_13_31_97), .A2(n_13_31_95), .A3(n_13_31_93), 
      .A4(n_13_31_92), .ZN(n_13_31_91));
   AOI22_X1 i_13_31_103 (.A1(\buffer[15][2][1] [10]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][1] [10]), .ZN(n_13_31_92));
   AOI22_X1 i_13_31_104 (.A1(\buffer[10][2][1] [10]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][1] [10]), .ZN(n_13_31_93));
   AOI22_X1 i_13_31_105 (.A1(\buffer[6][2][1] [10]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][1] [10]), .ZN(n_13_31_94));
   AOI22_X1 i_13_31_106 (.A1(\buffer[9][2][1] [10]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][1] [10]), .ZN(n_13_31_95));
   AOI22_X1 i_13_31_107 (.A1(\buffer[14][2][1] [10]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][1] [10]), .ZN(n_13_31_96));
   AOI22_X1 i_13_31_108 (.A1(\buffer[11][2][1] [10]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][1] [10]), .ZN(n_13_31_97));
   AOI22_X1 i_13_31_109 (.A1(\buffer[13][2][1] [10]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][1] [10]), .ZN(n_13_31_98));
   NAND4_X1 i_13_31_110 (.A1(n_13_31_107), .A2(n_13_31_105), .A3(n_13_31_103), 
      .A4(n_13_31_99), .ZN(\output_filter[2][1] [11]));
   AOI221_X1 i_13_31_111 (.A(n_13_31_100), .B1(n_25), .B2(\buffer[0][2][1] [11]), 
      .C1(\buffer[12][2][1] [11]), .C2(n_27), .ZN(n_13_31_99));
   NAND4_X1 i_13_31_112 (.A1(n_13_31_106), .A2(n_13_31_104), .A3(n_13_31_102), 
      .A4(n_13_31_101), .ZN(n_13_31_100));
   AOI22_X1 i_13_31_113 (.A1(\buffer[15][2][1] [11]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][1] [11]), .ZN(n_13_31_101));
   AOI22_X1 i_13_31_114 (.A1(\buffer[10][2][1] [11]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][1] [11]), .ZN(n_13_31_102));
   AOI22_X1 i_13_31_115 (.A1(\buffer[6][2][1] [11]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][1] [11]), .ZN(n_13_31_103));
   AOI22_X1 i_13_31_116 (.A1(\buffer[9][2][1] [11]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][2][1] [11]), .ZN(n_13_31_104));
   AOI22_X1 i_13_31_117 (.A1(\buffer[14][2][1] [11]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][1] [11]), .ZN(n_13_31_105));
   AOI22_X1 i_13_31_118 (.A1(\buffer[11][2][1] [11]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][1] [11]), .ZN(n_13_31_106));
   AOI22_X1 i_13_31_119 (.A1(\buffer[13][2][1] [11]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][2][1] [11]), .ZN(n_13_31_107));
   NAND4_X1 i_13_31_120 (.A1(n_13_31_116), .A2(n_13_31_114), .A3(n_13_31_112), 
      .A4(n_13_31_108), .ZN(\output_filter[2][1] [12]));
   AOI221_X1 i_13_31_121 (.A(n_13_31_109), .B1(n_25), .B2(\buffer[0][2][1] [12]), 
      .C1(\buffer[12][2][1] [12]), .C2(n_27), .ZN(n_13_31_108));
   NAND4_X1 i_13_31_122 (.A1(n_13_31_115), .A2(n_13_31_113), .A3(n_13_31_111), 
      .A4(n_13_31_110), .ZN(n_13_31_109));
   AOI22_X1 i_13_31_123 (.A1(\buffer[15][2][1] [12]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][1] [12]), .ZN(n_13_31_110));
   AOI22_X1 i_13_31_124 (.A1(\buffer[10][2][1] [12]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][1] [12]), .ZN(n_13_31_111));
   AOI22_X1 i_13_31_125 (.A1(\buffer[6][2][1] [12]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][1] [12]), .ZN(n_13_31_112));
   AOI22_X1 i_13_31_126 (.A1(\buffer[9][2][1] [12]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][1] [12]), .ZN(n_13_31_113));
   AOI22_X1 i_13_31_127 (.A1(\buffer[14][2][1] [12]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][1] [12]), .ZN(n_13_31_114));
   AOI22_X1 i_13_31_128 (.A1(\buffer[11][2][1] [12]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][1] [12]), .ZN(n_13_31_115));
   AOI22_X1 i_13_31_129 (.A1(\buffer[13][2][1] [12]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][1] [12]), .ZN(n_13_31_116));
   NAND4_X1 i_13_31_130 (.A1(n_13_31_125), .A2(n_13_31_123), .A3(n_13_31_121), 
      .A4(n_13_31_117), .ZN(\output_filter[2][1] [13]));
   AOI221_X1 i_13_31_131 (.A(n_13_31_118), .B1(n_25), .B2(\buffer[0][2][1] [13]), 
      .C1(\buffer[12][2][1] [13]), .C2(n_27), .ZN(n_13_31_117));
   NAND4_X1 i_13_31_132 (.A1(n_13_31_124), .A2(n_13_31_122), .A3(n_13_31_120), 
      .A4(n_13_31_119), .ZN(n_13_31_118));
   AOI22_X1 i_13_31_133 (.A1(\buffer[15][2][1] [13]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][1] [13]), .ZN(n_13_31_119));
   AOI22_X1 i_13_31_134 (.A1(\buffer[10][2][1] [13]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][1] [13]), .ZN(n_13_31_120));
   AOI22_X1 i_13_31_135 (.A1(\buffer[6][2][1] [13]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][1] [13]), .ZN(n_13_31_121));
   AOI22_X1 i_13_31_136 (.A1(\buffer[9][2][1] [13]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][2][1] [13]), .ZN(n_13_31_122));
   AOI22_X1 i_13_31_137 (.A1(\buffer[14][2][1] [13]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][1] [13]), .ZN(n_13_31_123));
   AOI22_X1 i_13_31_138 (.A1(\buffer[11][2][1] [13]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][1] [13]), .ZN(n_13_31_124));
   AOI22_X1 i_13_31_139 (.A1(\buffer[13][2][1] [13]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][2][1] [13]), .ZN(n_13_31_125));
   NAND4_X1 i_13_31_140 (.A1(n_13_31_134), .A2(n_13_31_132), .A3(n_13_31_130), 
      .A4(n_13_31_126), .ZN(\output_filter[2][1] [14]));
   AOI221_X1 i_13_31_141 (.A(n_13_31_127), .B1(n_25), .B2(\buffer[0][2][1] [14]), 
      .C1(\buffer[12][2][1] [14]), .C2(n_27), .ZN(n_13_31_126));
   NAND4_X1 i_13_31_142 (.A1(n_13_31_133), .A2(n_13_31_131), .A3(n_13_31_129), 
      .A4(n_13_31_128), .ZN(n_13_31_127));
   AOI22_X1 i_13_31_143 (.A1(\buffer[15][2][1] [14]), .A2(n_22), .B1(n_16), 
      .B2(\buffer[8][2][1] [14]), .ZN(n_13_31_128));
   AOI22_X1 i_13_31_144 (.A1(\buffer[10][2][1] [14]), .A2(n_21), .B1(n_29), 
      .B2(\buffer[7][2][1] [14]), .ZN(n_13_31_129));
   AOI22_X1 i_13_31_145 (.A1(\buffer[6][2][1] [14]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][1] [14]), .ZN(n_13_31_130));
   AOI22_X1 i_13_31_146 (.A1(\buffer[9][2][1] [14]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][1] [14]), .ZN(n_13_31_131));
   AOI22_X1 i_13_31_147 (.A1(\buffer[14][2][1] [14]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][1] [14]), .ZN(n_13_31_132));
   AOI22_X1 i_13_31_148 (.A1(\buffer[11][2][1] [14]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][1] [14]), .ZN(n_13_31_133));
   AOI22_X1 i_13_31_149 (.A1(\buffer[13][2][1] [14]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][1] [14]), .ZN(n_13_31_134));
   NAND2_X1 i_13_31_150 (.A1(n_13_31_137), .A2(n_13_31_135), .ZN(
      \output_filter[2][1] [15]));
   AOI221_X1 i_13_31_151 (.A(n_13_31_136), .B1(n_31), .B2(\buffer[3][2][1] [15]), 
      .C1(\buffer[14][2][1] [15]), .C2(n_19), .ZN(n_13_31_135));
   NAND3_X1 i_13_31_152 (.A1(n_13_31_143), .A2(n_13_31_141), .A3(n_13_31_139), 
      .ZN(n_13_31_136));
   AOI221_X1 i_13_31_153 (.A(n_13_31_138), .B1(n_16), .B2(\buffer[8][2][1] [15]), 
      .C1(\buffer[13][2][1] [15]), .C2(n_26), .ZN(n_13_31_137));
   NAND3_X1 i_13_31_154 (.A1(n_13_31_144), .A2(n_13_31_142), .A3(n_13_31_140), 
      .ZN(n_13_31_138));
   AOI22_X1 i_13_31_155 (.A1(\buffer[11][2][1] [15]), .A2(n_17), .B1(n_24), 
      .B2(\buffer[2][2][1] [15]), .ZN(n_13_31_139));
   AOI22_X1 i_13_31_156 (.A1(\buffer[10][2][1] [15]), .A2(n_21), .B1(n_23), 
      .B2(\buffer[1][2][1] [15]), .ZN(n_13_31_140));
   AOI22_X1 i_13_31_157 (.A1(\buffer[6][2][1] [15]), .A2(n_28), .B1(n_18), 
      .B2(\buffer[5][2][1] [15]), .ZN(n_13_31_141));
   AOI22_X1 i_13_31_158 (.A1(\buffer[9][2][1] [15]), .A2(n_20), .B1(n_30), 
      .B2(\buffer[4][2][1] [15]), .ZN(n_13_31_142));
   AOI22_X1 i_13_31_159 (.A1(\buffer[7][2][1] [15]), .A2(n_29), .B1(n_25), 
      .B2(\buffer[0][2][1] [15]), .ZN(n_13_31_143));
   AOI22_X1 i_13_31_160 (.A1(\buffer[15][2][1] [15]), .A2(n_22), .B1(n_27), 
      .B2(\buffer[12][2][1] [15]), .ZN(n_13_31_144));
   NAND4_X1 i_14_30_0 (.A1(n_14_30_8), .A2(n_14_30_6), .A3(n_14_30_4), .A4(
      n_14_30_0), .ZN(\output_filter[2][0] [0]));
   AOI221_X1 i_14_30_1 (.A(n_14_30_1), .B1(n_25), .B2(\buffer[0][2][0] [0]), 
      .C1(\buffer[12][2][0] [0]), .C2(n_27), .ZN(n_14_30_0));
   NAND4_X1 i_14_30_2 (.A1(n_14_30_7), .A2(n_14_30_5), .A3(n_14_30_3), .A4(
      n_14_30_2), .ZN(n_14_30_1));
   AOI22_X1 i_14_30_3 (.A1(\buffer[15][2][0] [0]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][0] [0]), .ZN(n_14_30_2));
   AOI22_X1 i_14_30_4 (.A1(\buffer[10][2][0] [0]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][0] [0]), .ZN(n_14_30_3));
   AOI22_X1 i_14_30_5 (.A1(\buffer[6][2][0] [0]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][2][0] [0]), .ZN(n_14_30_4));
   AOI22_X1 i_14_30_6 (.A1(\buffer[9][2][0] [0]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][2][0] [0]), .ZN(n_14_30_5));
   AOI22_X1 i_14_30_7 (.A1(\buffer[14][2][0] [0]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][0] [0]), .ZN(n_14_30_6));
   AOI22_X1 i_14_30_8 (.A1(\buffer[11][2][0] [0]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][0] [0]), .ZN(n_14_30_7));
   AOI22_X1 i_14_30_9 (.A1(\buffer[13][2][0] [0]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][0] [0]), .ZN(n_14_30_8));
   NAND4_X1 i_14_30_10 (.A1(n_14_30_17), .A2(n_14_30_15), .A3(n_14_30_13), 
      .A4(n_14_30_9), .ZN(\output_filter[2][0] [1]));
   AOI221_X1 i_14_30_11 (.A(n_14_30_10), .B1(n_25), .B2(\buffer[0][2][0] [1]), 
      .C1(\buffer[12][2][0] [1]), .C2(n_27), .ZN(n_14_30_9));
   NAND4_X1 i_14_30_12 (.A1(n_14_30_16), .A2(n_14_30_14), .A3(n_14_30_12), 
      .A4(n_14_30_11), .ZN(n_14_30_10));
   AOI22_X1 i_14_30_13 (.A1(\buffer[15][2][0] [1]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][0] [1]), .ZN(n_14_30_11));
   AOI22_X1 i_14_30_14 (.A1(\buffer[10][2][0] [1]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][0] [1]), .ZN(n_14_30_12));
   AOI22_X1 i_14_30_15 (.A1(\buffer[6][2][0] [1]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][0] [1]), .ZN(n_14_30_13));
   AOI22_X1 i_14_30_16 (.A1(\buffer[9][2][0] [1]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][0] [1]), .ZN(n_14_30_14));
   AOI22_X1 i_14_30_17 (.A1(\buffer[14][2][0] [1]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][0] [1]), .ZN(n_14_30_15));
   AOI22_X1 i_14_30_18 (.A1(\buffer[11][2][0] [1]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][0] [1]), .ZN(n_14_30_16));
   AOI22_X1 i_14_30_19 (.A1(\buffer[13][2][0] [1]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][0] [1]), .ZN(n_14_30_17));
   NAND4_X1 i_14_30_20 (.A1(n_14_30_26), .A2(n_14_30_24), .A3(n_14_30_22), 
      .A4(n_14_30_18), .ZN(\output_filter[2][0] [2]));
   AOI221_X1 i_14_30_21 (.A(n_14_30_19), .B1(n_25), .B2(\buffer[0][2][0] [2]), 
      .C1(\buffer[12][2][0] [2]), .C2(n_27), .ZN(n_14_30_18));
   NAND4_X1 i_14_30_22 (.A1(n_14_30_25), .A2(n_14_30_23), .A3(n_14_30_21), 
      .A4(n_14_30_20), .ZN(n_14_30_19));
   AOI22_X1 i_14_30_23 (.A1(\buffer[15][2][0] [2]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][0] [2]), .ZN(n_14_30_20));
   AOI22_X1 i_14_30_24 (.A1(\buffer[10][2][0] [2]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][0] [2]), .ZN(n_14_30_21));
   AOI22_X1 i_14_30_25 (.A1(\buffer[6][2][0] [2]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][0] [2]), .ZN(n_14_30_22));
   AOI22_X1 i_14_30_26 (.A1(\buffer[9][2][0] [2]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][0] [2]), .ZN(n_14_30_23));
   AOI22_X1 i_14_30_27 (.A1(\buffer[14][2][0] [2]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][0] [2]), .ZN(n_14_30_24));
   AOI22_X1 i_14_30_28 (.A1(\buffer[11][2][0] [2]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][0] [2]), .ZN(n_14_30_25));
   AOI22_X1 i_14_30_29 (.A1(\buffer[13][2][0] [2]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][0] [2]), .ZN(n_14_30_26));
   NAND4_X1 i_14_30_30 (.A1(n_14_30_35), .A2(n_14_30_33), .A3(n_14_30_31), 
      .A4(n_14_30_27), .ZN(\output_filter[2][0] [3]));
   AOI221_X1 i_14_30_31 (.A(n_14_30_28), .B1(n_25), .B2(\buffer[0][2][0] [3]), 
      .C1(\buffer[12][2][0] [3]), .C2(n_27), .ZN(n_14_30_27));
   NAND4_X1 i_14_30_32 (.A1(n_14_30_34), .A2(n_14_30_32), .A3(n_14_30_30), 
      .A4(n_14_30_29), .ZN(n_14_30_28));
   AOI22_X1 i_14_30_33 (.A1(\buffer[15][2][0] [3]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][0] [3]), .ZN(n_14_30_29));
   AOI22_X1 i_14_30_34 (.A1(\buffer[10][2][0] [3]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][0] [3]), .ZN(n_14_30_30));
   AOI22_X1 i_14_30_35 (.A1(\buffer[6][2][0] [3]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][0] [3]), .ZN(n_14_30_31));
   AOI22_X1 i_14_30_36 (.A1(\buffer[9][2][0] [3]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][0] [3]), .ZN(n_14_30_32));
   AOI22_X1 i_14_30_37 (.A1(\buffer[14][2][0] [3]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][0] [3]), .ZN(n_14_30_33));
   AOI22_X1 i_14_30_38 (.A1(\buffer[11][2][0] [3]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][0] [3]), .ZN(n_14_30_34));
   AOI22_X1 i_14_30_39 (.A1(\buffer[13][2][0] [3]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][0] [3]), .ZN(n_14_30_35));
   NAND4_X1 i_14_30_40 (.A1(n_14_30_44), .A2(n_14_30_42), .A3(n_14_30_40), 
      .A4(n_14_30_36), .ZN(\output_filter[2][0] [4]));
   AOI221_X1 i_14_30_41 (.A(n_14_30_37), .B1(n_25), .B2(\buffer[0][2][0] [4]), 
      .C1(\buffer[12][2][0] [4]), .C2(n_27), .ZN(n_14_30_36));
   NAND4_X1 i_14_30_42 (.A1(n_14_30_43), .A2(n_14_30_41), .A3(n_14_30_39), 
      .A4(n_14_30_38), .ZN(n_14_30_37));
   AOI22_X1 i_14_30_43 (.A1(\buffer[15][2][0] [4]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][0] [4]), .ZN(n_14_30_38));
   AOI22_X1 i_14_30_44 (.A1(\buffer[10][2][0] [4]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][0] [4]), .ZN(n_14_30_39));
   AOI22_X1 i_14_30_45 (.A1(\buffer[6][2][0] [4]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][0] [4]), .ZN(n_14_30_40));
   AOI22_X1 i_14_30_46 (.A1(\buffer[9][2][0] [4]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][2][0] [4]), .ZN(n_14_30_41));
   AOI22_X1 i_14_30_47 (.A1(\buffer[14][2][0] [4]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][0] [4]), .ZN(n_14_30_42));
   AOI22_X1 i_14_30_48 (.A1(\buffer[11][2][0] [4]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][0] [4]), .ZN(n_14_30_43));
   AOI22_X1 i_14_30_49 (.A1(\buffer[13][2][0] [4]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][2][0] [4]), .ZN(n_14_30_44));
   NAND4_X1 i_14_30_50 (.A1(n_14_30_53), .A2(n_14_30_51), .A3(n_14_30_49), 
      .A4(n_14_30_45), .ZN(\output_filter[2][0] [5]));
   AOI221_X1 i_14_30_51 (.A(n_14_30_46), .B1(n_25), .B2(\buffer[0][2][0] [5]), 
      .C1(\buffer[12][2][0] [5]), .C2(n_27), .ZN(n_14_30_45));
   NAND4_X1 i_14_30_52 (.A1(n_14_30_52), .A2(n_14_30_50), .A3(n_14_30_48), 
      .A4(n_14_30_47), .ZN(n_14_30_46));
   AOI22_X1 i_14_30_53 (.A1(\buffer[15][2][0] [5]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][0] [5]), .ZN(n_14_30_47));
   AOI22_X1 i_14_30_54 (.A1(\buffer[10][2][0] [5]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][0] [5]), .ZN(n_14_30_48));
   AOI22_X1 i_14_30_55 (.A1(\buffer[6][2][0] [5]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][0] [5]), .ZN(n_14_30_49));
   AOI22_X1 i_14_30_56 (.A1(\buffer[9][2][0] [5]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][0] [5]), .ZN(n_14_30_50));
   AOI22_X1 i_14_30_57 (.A1(\buffer[14][2][0] [5]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][0] [5]), .ZN(n_14_30_51));
   AOI22_X1 i_14_30_58 (.A1(\buffer[11][2][0] [5]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][0] [5]), .ZN(n_14_30_52));
   AOI22_X1 i_14_30_59 (.A1(\buffer[13][2][0] [5]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][0] [5]), .ZN(n_14_30_53));
   NAND4_X1 i_14_30_60 (.A1(n_14_30_62), .A2(n_14_30_60), .A3(n_14_30_58), 
      .A4(n_14_30_54), .ZN(\output_filter[2][0] [6]));
   AOI221_X1 i_14_30_61 (.A(n_14_30_55), .B1(n_25), .B2(\buffer[0][2][0] [6]), 
      .C1(\buffer[12][2][0] [6]), .C2(n_27), .ZN(n_14_30_54));
   NAND4_X1 i_14_30_62 (.A1(n_14_30_61), .A2(n_14_30_59), .A3(n_14_30_57), 
      .A4(n_14_30_56), .ZN(n_14_30_55));
   AOI22_X1 i_14_30_63 (.A1(\buffer[15][2][0] [6]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][0] [6]), .ZN(n_14_30_56));
   AOI22_X1 i_14_30_64 (.A1(\buffer[10][2][0] [6]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][0] [6]), .ZN(n_14_30_57));
   AOI22_X1 i_14_30_65 (.A1(\buffer[6][2][0] [6]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][0] [6]), .ZN(n_14_30_58));
   AOI22_X1 i_14_30_66 (.A1(\buffer[9][2][0] [6]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][0] [6]), .ZN(n_14_30_59));
   AOI22_X1 i_14_30_67 (.A1(\buffer[14][2][0] [6]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][0] [6]), .ZN(n_14_30_60));
   AOI22_X1 i_14_30_68 (.A1(\buffer[11][2][0] [6]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][0] [6]), .ZN(n_14_30_61));
   AOI22_X1 i_14_30_69 (.A1(\buffer[13][2][0] [6]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][0] [6]), .ZN(n_14_30_62));
   NAND4_X1 i_14_30_70 (.A1(n_14_30_71), .A2(n_14_30_69), .A3(n_14_30_67), 
      .A4(n_14_30_63), .ZN(\output_filter[2][0] [7]));
   AOI221_X1 i_14_30_71 (.A(n_14_30_64), .B1(n_25), .B2(\buffer[0][2][0] [7]), 
      .C1(\buffer[12][2][0] [7]), .C2(n_27), .ZN(n_14_30_63));
   NAND4_X1 i_14_30_72 (.A1(n_14_30_70), .A2(n_14_30_68), .A3(n_14_30_66), 
      .A4(n_14_30_65), .ZN(n_14_30_64));
   AOI22_X1 i_14_30_73 (.A1(\buffer[15][2][0] [7]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][0] [7]), .ZN(n_14_30_65));
   AOI22_X1 i_14_30_74 (.A1(\buffer[10][2][0] [7]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][0] [7]), .ZN(n_14_30_66));
   AOI22_X1 i_14_30_75 (.A1(\buffer[6][2][0] [7]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][0] [7]), .ZN(n_14_30_67));
   AOI22_X1 i_14_30_76 (.A1(\buffer[9][2][0] [7]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][2][0] [7]), .ZN(n_14_30_68));
   AOI22_X1 i_14_30_77 (.A1(\buffer[14][2][0] [7]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][0] [7]), .ZN(n_14_30_69));
   AOI22_X1 i_14_30_78 (.A1(\buffer[11][2][0] [7]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][0] [7]), .ZN(n_14_30_70));
   AOI22_X1 i_14_30_79 (.A1(\buffer[13][2][0] [7]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][2][0] [7]), .ZN(n_14_30_71));
   NAND4_X1 i_14_30_80 (.A1(n_14_30_80), .A2(n_14_30_78), .A3(n_14_30_76), 
      .A4(n_14_30_72), .ZN(\output_filter[2][0] [8]));
   AOI221_X1 i_14_30_81 (.A(n_14_30_73), .B1(n_25), .B2(\buffer[0][2][0] [8]), 
      .C1(\buffer[12][2][0] [8]), .C2(n_27), .ZN(n_14_30_72));
   NAND4_X1 i_14_30_82 (.A1(n_14_30_79), .A2(n_14_30_77), .A3(n_14_30_75), 
      .A4(n_14_30_74), .ZN(n_14_30_73));
   AOI22_X1 i_14_30_83 (.A1(\buffer[15][2][0] [8]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][0] [8]), .ZN(n_14_30_74));
   AOI22_X1 i_14_30_84 (.A1(\buffer[10][2][0] [8]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][0] [8]), .ZN(n_14_30_75));
   AOI22_X1 i_14_30_85 (.A1(\buffer[6][2][0] [8]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][0] [8]), .ZN(n_14_30_76));
   AOI22_X1 i_14_30_86 (.A1(\buffer[9][2][0] [8]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][0] [8]), .ZN(n_14_30_77));
   AOI22_X1 i_14_30_87 (.A1(\buffer[14][2][0] [8]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][0] [8]), .ZN(n_14_30_78));
   AOI22_X1 i_14_30_88 (.A1(\buffer[11][2][0] [8]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][0] [8]), .ZN(n_14_30_79));
   AOI22_X1 i_14_30_89 (.A1(\buffer[13][2][0] [8]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][0] [8]), .ZN(n_14_30_80));
   NAND4_X1 i_14_30_90 (.A1(n_14_30_89), .A2(n_14_30_87), .A3(n_14_30_85), 
      .A4(n_14_30_81), .ZN(\output_filter[2][0] [9]));
   AOI221_X1 i_14_30_91 (.A(n_14_30_82), .B1(n_25), .B2(\buffer[0][2][0] [9]), 
      .C1(\buffer[12][2][0] [9]), .C2(n_27), .ZN(n_14_30_81));
   NAND4_X1 i_14_30_92 (.A1(n_14_30_88), .A2(n_14_30_86), .A3(n_14_30_84), 
      .A4(n_14_30_83), .ZN(n_14_30_82));
   AOI22_X1 i_14_30_93 (.A1(\buffer[15][2][0] [9]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][0] [9]), .ZN(n_14_30_83));
   AOI22_X1 i_14_30_94 (.A1(\buffer[10][2][0] [9]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][0] [9]), .ZN(n_14_30_84));
   AOI22_X1 i_14_30_95 (.A1(\buffer[6][2][0] [9]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][0] [9]), .ZN(n_14_30_85));
   AOI22_X1 i_14_30_96 (.A1(\buffer[9][2][0] [9]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][2][0] [9]), .ZN(n_14_30_86));
   AOI22_X1 i_14_30_97 (.A1(\buffer[14][2][0] [9]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][0] [9]), .ZN(n_14_30_87));
   AOI22_X1 i_14_30_98 (.A1(\buffer[11][2][0] [9]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][0] [9]), .ZN(n_14_30_88));
   AOI22_X1 i_14_30_99 (.A1(\buffer[13][2][0] [9]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][2][0] [9]), .ZN(n_14_30_89));
   NAND4_X1 i_14_30_100 (.A1(n_14_30_98), .A2(n_14_30_96), .A3(n_14_30_94), 
      .A4(n_14_30_90), .ZN(\output_filter[2][0] [10]));
   AOI221_X1 i_14_30_101 (.A(n_14_30_91), .B1(n_25), .B2(\buffer[0][2][0] [10]), 
      .C1(\buffer[12][2][0] [10]), .C2(n_27), .ZN(n_14_30_90));
   NAND4_X1 i_14_30_102 (.A1(n_14_30_97), .A2(n_14_30_95), .A3(n_14_30_93), 
      .A4(n_14_30_92), .ZN(n_14_30_91));
   AOI22_X1 i_14_30_103 (.A1(\buffer[15][2][0] [10]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][0] [10]), .ZN(n_14_30_92));
   AOI22_X1 i_14_30_104 (.A1(\buffer[10][2][0] [10]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][0] [10]), .ZN(n_14_30_93));
   AOI22_X1 i_14_30_105 (.A1(\buffer[6][2][0] [10]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][0] [10]), .ZN(n_14_30_94));
   AOI22_X1 i_14_30_106 (.A1(\buffer[9][2][0] [10]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][0] [10]), .ZN(n_14_30_95));
   AOI22_X1 i_14_30_107 (.A1(\buffer[14][2][0] [10]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][0] [10]), .ZN(n_14_30_96));
   AOI22_X1 i_14_30_108 (.A1(\buffer[11][2][0] [10]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][0] [10]), .ZN(n_14_30_97));
   AOI22_X1 i_14_30_109 (.A1(\buffer[13][2][0] [10]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][0] [10]), .ZN(n_14_30_98));
   NAND4_X1 i_14_30_110 (.A1(n_14_30_107), .A2(n_14_30_105), .A3(n_14_30_103), 
      .A4(n_14_30_99), .ZN(\output_filter[2][0] [11]));
   AOI221_X1 i_14_30_111 (.A(n_14_30_100), .B1(n_25), .B2(\buffer[0][2][0] [11]), 
      .C1(\buffer[12][2][0] [11]), .C2(n_27), .ZN(n_14_30_99));
   NAND4_X1 i_14_30_112 (.A1(n_14_30_106), .A2(n_14_30_104), .A3(n_14_30_102), 
      .A4(n_14_30_101), .ZN(n_14_30_100));
   AOI22_X1 i_14_30_113 (.A1(\buffer[15][2][0] [11]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][0] [11]), .ZN(n_14_30_101));
   AOI22_X1 i_14_30_114 (.A1(\buffer[10][2][0] [11]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][0] [11]), .ZN(n_14_30_102));
   AOI22_X1 i_14_30_115 (.A1(\buffer[6][2][0] [11]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][0] [11]), .ZN(n_14_30_103));
   AOI22_X1 i_14_30_116 (.A1(\buffer[9][2][0] [11]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][2][0] [11]), .ZN(n_14_30_104));
   AOI22_X1 i_14_30_117 (.A1(\buffer[14][2][0] [11]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][0] [11]), .ZN(n_14_30_105));
   AOI22_X1 i_14_30_118 (.A1(\buffer[11][2][0] [11]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][0] [11]), .ZN(n_14_30_106));
   AOI22_X1 i_14_30_119 (.A1(\buffer[13][2][0] [11]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][2][0] [11]), .ZN(n_14_30_107));
   NAND4_X1 i_14_30_120 (.A1(n_14_30_116), .A2(n_14_30_114), .A3(n_14_30_112), 
      .A4(n_14_30_108), .ZN(\output_filter[2][0] [12]));
   AOI221_X1 i_14_30_121 (.A(n_14_30_109), .B1(n_25), .B2(\buffer[0][2][0] [12]), 
      .C1(\buffer[12][2][0] [12]), .C2(n_27), .ZN(n_14_30_108));
   NAND4_X1 i_14_30_122 (.A1(n_14_30_115), .A2(n_14_30_113), .A3(n_14_30_111), 
      .A4(n_14_30_110), .ZN(n_14_30_109));
   AOI22_X1 i_14_30_123 (.A1(\buffer[15][2][0] [12]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][0] [12]), .ZN(n_14_30_110));
   AOI22_X1 i_14_30_124 (.A1(\buffer[10][2][0] [12]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][0] [12]), .ZN(n_14_30_111));
   AOI22_X1 i_14_30_125 (.A1(\buffer[6][2][0] [12]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][0] [12]), .ZN(n_14_30_112));
   AOI22_X1 i_14_30_126 (.A1(\buffer[9][2][0] [12]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][0] [12]), .ZN(n_14_30_113));
   AOI22_X1 i_14_30_127 (.A1(\buffer[14][2][0] [12]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][0] [12]), .ZN(n_14_30_114));
   AOI22_X1 i_14_30_128 (.A1(\buffer[11][2][0] [12]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][0] [12]), .ZN(n_14_30_115));
   AOI22_X1 i_14_30_129 (.A1(\buffer[13][2][0] [12]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][0] [12]), .ZN(n_14_30_116));
   NAND4_X1 i_14_30_130 (.A1(n_14_30_125), .A2(n_14_30_123), .A3(n_14_30_121), 
      .A4(n_14_30_117), .ZN(\output_filter[2][0] [13]));
   AOI221_X1 i_14_30_131 (.A(n_14_30_118), .B1(n_25), .B2(\buffer[0][2][0] [13]), 
      .C1(\buffer[12][2][0] [13]), .C2(n_27), .ZN(n_14_30_117));
   NAND4_X1 i_14_30_132 (.A1(n_14_30_124), .A2(n_14_30_122), .A3(n_14_30_120), 
      .A4(n_14_30_119), .ZN(n_14_30_118));
   AOI22_X1 i_14_30_133 (.A1(\buffer[15][2][0] [13]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][0] [13]), .ZN(n_14_30_119));
   AOI22_X1 i_14_30_134 (.A1(\buffer[10][2][0] [13]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][0] [13]), .ZN(n_14_30_120));
   AOI22_X1 i_14_30_135 (.A1(\buffer[6][2][0] [13]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][0] [13]), .ZN(n_14_30_121));
   AOI22_X1 i_14_30_136 (.A1(\buffer[9][2][0] [13]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][2][0] [13]), .ZN(n_14_30_122));
   AOI22_X1 i_14_30_137 (.A1(\buffer[14][2][0] [13]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][0] [13]), .ZN(n_14_30_123));
   AOI22_X1 i_14_30_138 (.A1(\buffer[11][2][0] [13]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][0] [13]), .ZN(n_14_30_124));
   AOI22_X1 i_14_30_139 (.A1(\buffer[13][2][0] [13]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][2][0] [13]), .ZN(n_14_30_125));
   NAND4_X1 i_14_30_140 (.A1(n_14_30_134), .A2(n_14_30_132), .A3(n_14_30_130), 
      .A4(n_14_30_126), .ZN(\output_filter[2][0] [14]));
   AOI221_X1 i_14_30_141 (.A(n_14_30_127), .B1(n_25), .B2(\buffer[0][2][0] [14]), 
      .C1(\buffer[12][2][0] [14]), .C2(n_27), .ZN(n_14_30_126));
   NAND4_X1 i_14_30_142 (.A1(n_14_30_133), .A2(n_14_30_131), .A3(n_14_30_129), 
      .A4(n_14_30_128), .ZN(n_14_30_127));
   AOI22_X1 i_14_30_143 (.A1(\buffer[15][2][0] [14]), .A2(n_22), .B1(n_16), 
      .B2(\buffer[8][2][0] [14]), .ZN(n_14_30_128));
   AOI22_X1 i_14_30_144 (.A1(\buffer[10][2][0] [14]), .A2(n_21), .B1(n_29), 
      .B2(\buffer[7][2][0] [14]), .ZN(n_14_30_129));
   AOI22_X1 i_14_30_145 (.A1(\buffer[6][2][0] [14]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][0] [14]), .ZN(n_14_30_130));
   AOI22_X1 i_14_30_146 (.A1(\buffer[9][2][0] [14]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][0] [14]), .ZN(n_14_30_131));
   AOI22_X1 i_14_30_147 (.A1(\buffer[14][2][0] [14]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][0] [14]), .ZN(n_14_30_132));
   AOI22_X1 i_14_30_148 (.A1(\buffer[11][2][0] [14]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][0] [14]), .ZN(n_14_30_133));
   AOI22_X1 i_14_30_149 (.A1(\buffer[13][2][0] [14]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][0] [14]), .ZN(n_14_30_134));
   NAND2_X1 i_14_30_150 (.A1(n_14_30_137), .A2(n_14_30_135), .ZN(
      \output_filter[2][0] [15]));
   AOI221_X1 i_14_30_151 (.A(n_14_30_136), .B1(n_31), .B2(\buffer[3][2][0] [15]), 
      .C1(\buffer[14][2][0] [15]), .C2(n_19), .ZN(n_14_30_135));
   NAND3_X1 i_14_30_152 (.A1(n_14_30_143), .A2(n_14_30_141), .A3(n_14_30_139), 
      .ZN(n_14_30_136));
   AOI221_X1 i_14_30_153 (.A(n_14_30_138), .B1(n_16), .B2(\buffer[8][2][0] [15]), 
      .C1(\buffer[13][2][0] [15]), .C2(n_26), .ZN(n_14_30_137));
   NAND3_X1 i_14_30_154 (.A1(n_14_30_144), .A2(n_14_30_142), .A3(n_14_30_140), 
      .ZN(n_14_30_138));
   AOI22_X1 i_14_30_155 (.A1(\buffer[11][2][0] [15]), .A2(n_17), .B1(n_24), 
      .B2(\buffer[2][2][0] [15]), .ZN(n_14_30_139));
   AOI22_X1 i_14_30_156 (.A1(\buffer[10][2][0] [15]), .A2(n_21), .B1(n_23), 
      .B2(\buffer[1][2][0] [15]), .ZN(n_14_30_140));
   AOI22_X1 i_14_30_157 (.A1(\buffer[6][2][0] [15]), .A2(n_28), .B1(n_18), 
      .B2(\buffer[5][2][0] [15]), .ZN(n_14_30_141));
   AOI22_X1 i_14_30_158 (.A1(\buffer[9][2][0] [15]), .A2(n_20), .B1(n_30), 
      .B2(\buffer[4][2][0] [15]), .ZN(n_14_30_142));
   AOI22_X1 i_14_30_159 (.A1(\buffer[7][2][0] [15]), .A2(n_29), .B1(n_25), 
      .B2(\buffer[0][2][0] [15]), .ZN(n_14_30_143));
   AOI22_X1 i_14_30_160 (.A1(\buffer[15][2][0] [15]), .A2(n_22), .B1(n_27), 
      .B2(\buffer[12][2][0] [15]), .ZN(n_14_30_144));
   NAND4_X1 i_15_29_0 (.A1(n_15_29_8), .A2(n_15_29_6), .A3(n_15_29_4), .A4(
      n_15_29_0), .ZN(\output_filter[1][4] [0]));
   AOI221_X1 i_15_29_1 (.A(n_15_29_1), .B1(n_25), .B2(\buffer[0][1][4] [0]), 
      .C1(\buffer[12][1][4] [0]), .C2(n_27), .ZN(n_15_29_0));
   NAND4_X1 i_15_29_2 (.A1(n_15_29_7), .A2(n_15_29_5), .A3(n_15_29_3), .A4(
      n_15_29_2), .ZN(n_15_29_1));
   AOI22_X1 i_15_29_3 (.A1(\buffer[15][1][4] [0]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][4] [0]), .ZN(n_15_29_2));
   AOI22_X1 i_15_29_4 (.A1(\buffer[10][1][4] [0]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][4] [0]), .ZN(n_15_29_3));
   AOI22_X1 i_15_29_5 (.A1(\buffer[6][1][4] [0]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][1][4] [0]), .ZN(n_15_29_4));
   AOI22_X1 i_15_29_6 (.A1(\buffer[9][1][4] [0]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][1][4] [0]), .ZN(n_15_29_5));
   AOI22_X1 i_15_29_7 (.A1(\buffer[14][1][4] [0]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][4] [0]), .ZN(n_15_29_6));
   AOI22_X1 i_15_29_8 (.A1(\buffer[11][1][4] [0]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][4] [0]), .ZN(n_15_29_7));
   AOI22_X1 i_15_29_9 (.A1(\buffer[13][1][4] [0]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][4] [0]), .ZN(n_15_29_8));
   NAND4_X1 i_15_29_10 (.A1(n_15_29_17), .A2(n_15_29_15), .A3(n_15_29_13), 
      .A4(n_15_29_9), .ZN(\output_filter[1][4] [1]));
   AOI221_X1 i_15_29_11 (.A(n_15_29_10), .B1(n_25), .B2(\buffer[0][1][4] [1]), 
      .C1(\buffer[12][1][4] [1]), .C2(n_27), .ZN(n_15_29_9));
   NAND4_X1 i_15_29_12 (.A1(n_15_29_16), .A2(n_15_29_14), .A3(n_15_29_12), 
      .A4(n_15_29_11), .ZN(n_15_29_10));
   AOI22_X1 i_15_29_13 (.A1(\buffer[15][1][4] [1]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][4] [1]), .ZN(n_15_29_11));
   AOI22_X1 i_15_29_14 (.A1(\buffer[10][1][4] [1]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][4] [1]), .ZN(n_15_29_12));
   AOI22_X1 i_15_29_15 (.A1(\buffer[6][1][4] [1]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][4] [1]), .ZN(n_15_29_13));
   AOI22_X1 i_15_29_16 (.A1(\buffer[9][1][4] [1]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][4] [1]), .ZN(n_15_29_14));
   AOI22_X1 i_15_29_17 (.A1(\buffer[14][1][4] [1]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][4] [1]), .ZN(n_15_29_15));
   AOI22_X1 i_15_29_18 (.A1(\buffer[11][1][4] [1]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][4] [1]), .ZN(n_15_29_16));
   AOI22_X1 i_15_29_19 (.A1(\buffer[13][1][4] [1]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][4] [1]), .ZN(n_15_29_17));
   NAND4_X1 i_15_29_20 (.A1(n_15_29_26), .A2(n_15_29_24), .A3(n_15_29_22), 
      .A4(n_15_29_18), .ZN(\output_filter[1][4] [2]));
   AOI221_X1 i_15_29_21 (.A(n_15_29_19), .B1(n_25), .B2(\buffer[0][1][4] [2]), 
      .C1(\buffer[12][1][4] [2]), .C2(n_27), .ZN(n_15_29_18));
   NAND4_X1 i_15_29_22 (.A1(n_15_29_25), .A2(n_15_29_23), .A3(n_15_29_21), 
      .A4(n_15_29_20), .ZN(n_15_29_19));
   AOI22_X1 i_15_29_23 (.A1(\buffer[15][1][4] [2]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][4] [2]), .ZN(n_15_29_20));
   AOI22_X1 i_15_29_24 (.A1(\buffer[10][1][4] [2]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][4] [2]), .ZN(n_15_29_21));
   AOI22_X1 i_15_29_25 (.A1(\buffer[6][1][4] [2]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][4] [2]), .ZN(n_15_29_22));
   AOI22_X1 i_15_29_26 (.A1(\buffer[9][1][4] [2]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][4] [2]), .ZN(n_15_29_23));
   AOI22_X1 i_15_29_27 (.A1(\buffer[14][1][4] [2]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][4] [2]), .ZN(n_15_29_24));
   AOI22_X1 i_15_29_28 (.A1(\buffer[11][1][4] [2]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][4] [2]), .ZN(n_15_29_25));
   AOI22_X1 i_15_29_29 (.A1(\buffer[13][1][4] [2]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][4] [2]), .ZN(n_15_29_26));
   NAND4_X1 i_15_29_30 (.A1(n_15_29_35), .A2(n_15_29_33), .A3(n_15_29_31), 
      .A4(n_15_29_27), .ZN(\output_filter[1][4] [3]));
   AOI221_X1 i_15_29_31 (.A(n_15_29_28), .B1(n_25), .B2(\buffer[0][1][4] [3]), 
      .C1(\buffer[12][1][4] [3]), .C2(n_27), .ZN(n_15_29_27));
   NAND4_X1 i_15_29_32 (.A1(n_15_29_34), .A2(n_15_29_32), .A3(n_15_29_30), 
      .A4(n_15_29_29), .ZN(n_15_29_28));
   AOI22_X1 i_15_29_33 (.A1(\buffer[15][1][4] [3]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][4] [3]), .ZN(n_15_29_29));
   AOI22_X1 i_15_29_34 (.A1(\buffer[10][1][4] [3]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][4] [3]), .ZN(n_15_29_30));
   AOI22_X1 i_15_29_35 (.A1(\buffer[6][1][4] [3]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][4] [3]), .ZN(n_15_29_31));
   AOI22_X1 i_15_29_36 (.A1(\buffer[9][1][4] [3]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][4] [3]), .ZN(n_15_29_32));
   AOI22_X1 i_15_29_37 (.A1(\buffer[14][1][4] [3]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][4] [3]), .ZN(n_15_29_33));
   AOI22_X1 i_15_29_38 (.A1(\buffer[11][1][4] [3]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][4] [3]), .ZN(n_15_29_34));
   AOI22_X1 i_15_29_39 (.A1(\buffer[13][1][4] [3]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][4] [3]), .ZN(n_15_29_35));
   NAND4_X1 i_15_29_40 (.A1(n_15_29_44), .A2(n_15_29_42), .A3(n_15_29_40), 
      .A4(n_15_29_36), .ZN(\output_filter[1][4] [4]));
   AOI221_X1 i_15_29_41 (.A(n_15_29_37), .B1(n_25), .B2(\buffer[0][1][4] [4]), 
      .C1(\buffer[12][1][4] [4]), .C2(n_27), .ZN(n_15_29_36));
   NAND4_X1 i_15_29_42 (.A1(n_15_29_43), .A2(n_15_29_41), .A3(n_15_29_39), 
      .A4(n_15_29_38), .ZN(n_15_29_37));
   AOI22_X1 i_15_29_43 (.A1(\buffer[15][1][4] [4]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][4] [4]), .ZN(n_15_29_38));
   AOI22_X1 i_15_29_44 (.A1(\buffer[10][1][4] [4]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][4] [4]), .ZN(n_15_29_39));
   AOI22_X1 i_15_29_45 (.A1(\buffer[6][1][4] [4]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][4] [4]), .ZN(n_15_29_40));
   AOI22_X1 i_15_29_46 (.A1(\buffer[9][1][4] [4]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][1][4] [4]), .ZN(n_15_29_41));
   AOI22_X1 i_15_29_47 (.A1(\buffer[14][1][4] [4]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][4] [4]), .ZN(n_15_29_42));
   AOI22_X1 i_15_29_48 (.A1(\buffer[11][1][4] [4]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][4] [4]), .ZN(n_15_29_43));
   AOI22_X1 i_15_29_49 (.A1(\buffer[13][1][4] [4]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][1][4] [4]), .ZN(n_15_29_44));
   NAND4_X1 i_15_29_50 (.A1(n_15_29_53), .A2(n_15_29_51), .A3(n_15_29_49), 
      .A4(n_15_29_45), .ZN(\output_filter[1][4] [5]));
   AOI221_X1 i_15_29_51 (.A(n_15_29_46), .B1(n_25), .B2(\buffer[0][1][4] [5]), 
      .C1(\buffer[12][1][4] [5]), .C2(n_27), .ZN(n_15_29_45));
   NAND4_X1 i_15_29_52 (.A1(n_15_29_52), .A2(n_15_29_50), .A3(n_15_29_48), 
      .A4(n_15_29_47), .ZN(n_15_29_46));
   AOI22_X1 i_15_29_53 (.A1(\buffer[15][1][4] [5]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][4] [5]), .ZN(n_15_29_47));
   AOI22_X1 i_15_29_54 (.A1(\buffer[10][1][4] [5]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][4] [5]), .ZN(n_15_29_48));
   AOI22_X1 i_15_29_55 (.A1(\buffer[6][1][4] [5]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][4] [5]), .ZN(n_15_29_49));
   AOI22_X1 i_15_29_56 (.A1(\buffer[9][1][4] [5]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][4] [5]), .ZN(n_15_29_50));
   AOI22_X1 i_15_29_57 (.A1(\buffer[14][1][4] [5]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][4] [5]), .ZN(n_15_29_51));
   AOI22_X1 i_15_29_58 (.A1(\buffer[11][1][4] [5]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][4] [5]), .ZN(n_15_29_52));
   AOI22_X1 i_15_29_59 (.A1(\buffer[13][1][4] [5]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][4] [5]), .ZN(n_15_29_53));
   NAND4_X1 i_15_29_60 (.A1(n_15_29_62), .A2(n_15_29_60), .A3(n_15_29_58), 
      .A4(n_15_29_54), .ZN(\output_filter[1][4] [6]));
   AOI221_X1 i_15_29_61 (.A(n_15_29_55), .B1(n_25), .B2(\buffer[0][1][4] [6]), 
      .C1(\buffer[12][1][4] [6]), .C2(n_27), .ZN(n_15_29_54));
   NAND4_X1 i_15_29_62 (.A1(n_15_29_61), .A2(n_15_29_59), .A3(n_15_29_57), 
      .A4(n_15_29_56), .ZN(n_15_29_55));
   AOI22_X1 i_15_29_63 (.A1(\buffer[15][1][4] [6]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][4] [6]), .ZN(n_15_29_56));
   AOI22_X1 i_15_29_64 (.A1(\buffer[10][1][4] [6]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][4] [6]), .ZN(n_15_29_57));
   AOI22_X1 i_15_29_65 (.A1(\buffer[6][1][4] [6]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][4] [6]), .ZN(n_15_29_58));
   AOI22_X1 i_15_29_66 (.A1(\buffer[9][1][4] [6]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][4] [6]), .ZN(n_15_29_59));
   AOI22_X1 i_15_29_67 (.A1(\buffer[14][1][4] [6]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][4] [6]), .ZN(n_15_29_60));
   AOI22_X1 i_15_29_68 (.A1(\buffer[11][1][4] [6]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][4] [6]), .ZN(n_15_29_61));
   AOI22_X1 i_15_29_69 (.A1(\buffer[13][1][4] [6]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][4] [6]), .ZN(n_15_29_62));
   NAND4_X1 i_15_29_70 (.A1(n_15_29_71), .A2(n_15_29_69), .A3(n_15_29_67), 
      .A4(n_15_29_63), .ZN(\output_filter[1][4] [7]));
   AOI221_X1 i_15_29_71 (.A(n_15_29_64), .B1(n_25), .B2(\buffer[0][1][4] [7]), 
      .C1(\buffer[12][1][4] [7]), .C2(n_27), .ZN(n_15_29_63));
   NAND4_X1 i_15_29_72 (.A1(n_15_29_70), .A2(n_15_29_68), .A3(n_15_29_66), 
      .A4(n_15_29_65), .ZN(n_15_29_64));
   AOI22_X1 i_15_29_73 (.A1(\buffer[15][1][4] [7]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][4] [7]), .ZN(n_15_29_65));
   AOI22_X1 i_15_29_74 (.A1(\buffer[10][1][4] [7]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][4] [7]), .ZN(n_15_29_66));
   AOI22_X1 i_15_29_75 (.A1(\buffer[6][1][4] [7]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][4] [7]), .ZN(n_15_29_67));
   AOI22_X1 i_15_29_76 (.A1(\buffer[9][1][4] [7]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][1][4] [7]), .ZN(n_15_29_68));
   AOI22_X1 i_15_29_77 (.A1(\buffer[14][1][4] [7]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][4] [7]), .ZN(n_15_29_69));
   AOI22_X1 i_15_29_78 (.A1(\buffer[11][1][4] [7]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][4] [7]), .ZN(n_15_29_70));
   AOI22_X1 i_15_29_79 (.A1(\buffer[13][1][4] [7]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][1][4] [7]), .ZN(n_15_29_71));
   NAND4_X1 i_15_29_80 (.A1(n_15_29_80), .A2(n_15_29_78), .A3(n_15_29_76), 
      .A4(n_15_29_72), .ZN(\output_filter[1][4] [8]));
   AOI221_X1 i_15_29_81 (.A(n_15_29_73), .B1(n_25), .B2(\buffer[0][1][4] [8]), 
      .C1(\buffer[12][1][4] [8]), .C2(n_27), .ZN(n_15_29_72));
   NAND4_X1 i_15_29_82 (.A1(n_15_29_79), .A2(n_15_29_77), .A3(n_15_29_75), 
      .A4(n_15_29_74), .ZN(n_15_29_73));
   AOI22_X1 i_15_29_83 (.A1(\buffer[15][1][4] [8]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][4] [8]), .ZN(n_15_29_74));
   AOI22_X1 i_15_29_84 (.A1(\buffer[10][1][4] [8]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][4] [8]), .ZN(n_15_29_75));
   AOI22_X1 i_15_29_85 (.A1(\buffer[6][1][4] [8]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][4] [8]), .ZN(n_15_29_76));
   AOI22_X1 i_15_29_86 (.A1(\buffer[9][1][4] [8]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][4] [8]), .ZN(n_15_29_77));
   AOI22_X1 i_15_29_87 (.A1(\buffer[14][1][4] [8]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][4] [8]), .ZN(n_15_29_78));
   AOI22_X1 i_15_29_88 (.A1(\buffer[11][1][4] [8]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][4] [8]), .ZN(n_15_29_79));
   AOI22_X1 i_15_29_89 (.A1(\buffer[13][1][4] [8]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][4] [8]), .ZN(n_15_29_80));
   NAND4_X1 i_15_29_90 (.A1(n_15_29_89), .A2(n_15_29_87), .A3(n_15_29_85), 
      .A4(n_15_29_81), .ZN(\output_filter[1][4] [9]));
   AOI221_X1 i_15_29_91 (.A(n_15_29_82), .B1(n_25), .B2(\buffer[0][1][4] [9]), 
      .C1(\buffer[12][1][4] [9]), .C2(n_27), .ZN(n_15_29_81));
   NAND4_X1 i_15_29_92 (.A1(n_15_29_88), .A2(n_15_29_86), .A3(n_15_29_84), 
      .A4(n_15_29_83), .ZN(n_15_29_82));
   AOI22_X1 i_15_29_93 (.A1(\buffer[15][1][4] [9]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][4] [9]), .ZN(n_15_29_83));
   AOI22_X1 i_15_29_94 (.A1(\buffer[10][1][4] [9]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][4] [9]), .ZN(n_15_29_84));
   AOI22_X1 i_15_29_95 (.A1(\buffer[6][1][4] [9]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][4] [9]), .ZN(n_15_29_85));
   AOI22_X1 i_15_29_96 (.A1(\buffer[9][1][4] [9]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][1][4] [9]), .ZN(n_15_29_86));
   AOI22_X1 i_15_29_97 (.A1(\buffer[14][1][4] [9]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][4] [9]), .ZN(n_15_29_87));
   AOI22_X1 i_15_29_98 (.A1(\buffer[11][1][4] [9]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][4] [9]), .ZN(n_15_29_88));
   AOI22_X1 i_15_29_99 (.A1(\buffer[13][1][4] [9]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][1][4] [9]), .ZN(n_15_29_89));
   NAND4_X1 i_15_29_100 (.A1(n_15_29_98), .A2(n_15_29_96), .A3(n_15_29_94), 
      .A4(n_15_29_90), .ZN(\output_filter[1][4] [10]));
   AOI221_X1 i_15_29_101 (.A(n_15_29_91), .B1(n_25), .B2(\buffer[0][1][4] [10]), 
      .C1(\buffer[12][1][4] [10]), .C2(n_27), .ZN(n_15_29_90));
   NAND4_X1 i_15_29_102 (.A1(n_15_29_97), .A2(n_15_29_95), .A3(n_15_29_93), 
      .A4(n_15_29_92), .ZN(n_15_29_91));
   AOI22_X1 i_15_29_103 (.A1(\buffer[15][1][4] [10]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][4] [10]), .ZN(n_15_29_92));
   AOI22_X1 i_15_29_104 (.A1(\buffer[10][1][4] [10]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][4] [10]), .ZN(n_15_29_93));
   AOI22_X1 i_15_29_105 (.A1(\buffer[6][1][4] [10]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][4] [10]), .ZN(n_15_29_94));
   AOI22_X1 i_15_29_106 (.A1(\buffer[9][1][4] [10]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][4] [10]), .ZN(n_15_29_95));
   AOI22_X1 i_15_29_107 (.A1(\buffer[14][1][4] [10]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][4] [10]), .ZN(n_15_29_96));
   AOI22_X1 i_15_29_108 (.A1(\buffer[11][1][4] [10]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][4] [10]), .ZN(n_15_29_97));
   AOI22_X1 i_15_29_109 (.A1(\buffer[13][1][4] [10]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][4] [10]), .ZN(n_15_29_98));
   NAND4_X1 i_15_29_110 (.A1(n_15_29_107), .A2(n_15_29_105), .A3(n_15_29_103), 
      .A4(n_15_29_99), .ZN(\output_filter[1][4] [11]));
   AOI221_X1 i_15_29_111 (.A(n_15_29_100), .B1(n_25), .B2(\buffer[0][1][4] [11]), 
      .C1(\buffer[12][1][4] [11]), .C2(n_27), .ZN(n_15_29_99));
   NAND4_X1 i_15_29_112 (.A1(n_15_29_106), .A2(n_15_29_104), .A3(n_15_29_102), 
      .A4(n_15_29_101), .ZN(n_15_29_100));
   AOI22_X1 i_15_29_113 (.A1(\buffer[15][1][4] [11]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][4] [11]), .ZN(n_15_29_101));
   AOI22_X1 i_15_29_114 (.A1(\buffer[10][1][4] [11]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][4] [11]), .ZN(n_15_29_102));
   AOI22_X1 i_15_29_115 (.A1(\buffer[6][1][4] [11]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][4] [11]), .ZN(n_15_29_103));
   AOI22_X1 i_15_29_116 (.A1(\buffer[9][1][4] [11]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][1][4] [11]), .ZN(n_15_29_104));
   AOI22_X1 i_15_29_117 (.A1(\buffer[14][1][4] [11]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][4] [11]), .ZN(n_15_29_105));
   AOI22_X1 i_15_29_118 (.A1(\buffer[11][1][4] [11]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][4] [11]), .ZN(n_15_29_106));
   AOI22_X1 i_15_29_119 (.A1(\buffer[13][1][4] [11]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][1][4] [11]), .ZN(n_15_29_107));
   NAND4_X1 i_15_29_120 (.A1(n_15_29_116), .A2(n_15_29_114), .A3(n_15_29_112), 
      .A4(n_15_29_108), .ZN(\output_filter[1][4] [12]));
   AOI221_X1 i_15_29_121 (.A(n_15_29_109), .B1(n_25), .B2(\buffer[0][1][4] [12]), 
      .C1(\buffer[12][1][4] [12]), .C2(n_27), .ZN(n_15_29_108));
   NAND4_X1 i_15_29_122 (.A1(n_15_29_115), .A2(n_15_29_113), .A3(n_15_29_111), 
      .A4(n_15_29_110), .ZN(n_15_29_109));
   AOI22_X1 i_15_29_123 (.A1(\buffer[15][1][4] [12]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][4] [12]), .ZN(n_15_29_110));
   AOI22_X1 i_15_29_124 (.A1(\buffer[10][1][4] [12]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][4] [12]), .ZN(n_15_29_111));
   AOI22_X1 i_15_29_125 (.A1(\buffer[6][1][4] [12]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][4] [12]), .ZN(n_15_29_112));
   AOI22_X1 i_15_29_126 (.A1(\buffer[9][1][4] [12]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][4] [12]), .ZN(n_15_29_113));
   AOI22_X1 i_15_29_127 (.A1(\buffer[14][1][4] [12]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][4] [12]), .ZN(n_15_29_114));
   AOI22_X1 i_15_29_128 (.A1(\buffer[11][1][4] [12]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][4] [12]), .ZN(n_15_29_115));
   AOI22_X1 i_15_29_129 (.A1(\buffer[13][1][4] [12]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][4] [12]), .ZN(n_15_29_116));
   NAND4_X1 i_15_29_130 (.A1(n_15_29_125), .A2(n_15_29_123), .A3(n_15_29_121), 
      .A4(n_15_29_117), .ZN(\output_filter[1][4] [13]));
   AOI221_X1 i_15_29_131 (.A(n_15_29_118), .B1(n_25), .B2(\buffer[0][1][4] [13]), 
      .C1(\buffer[12][1][4] [13]), .C2(n_27), .ZN(n_15_29_117));
   NAND4_X1 i_15_29_132 (.A1(n_15_29_124), .A2(n_15_29_122), .A3(n_15_29_120), 
      .A4(n_15_29_119), .ZN(n_15_29_118));
   AOI22_X1 i_15_29_133 (.A1(\buffer[15][1][4] [13]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][4] [13]), .ZN(n_15_29_119));
   AOI22_X1 i_15_29_134 (.A1(\buffer[10][1][4] [13]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][4] [13]), .ZN(n_15_29_120));
   AOI22_X1 i_15_29_135 (.A1(\buffer[6][1][4] [13]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][4] [13]), .ZN(n_15_29_121));
   AOI22_X1 i_15_29_136 (.A1(\buffer[9][1][4] [13]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][1][4] [13]), .ZN(n_15_29_122));
   AOI22_X1 i_15_29_137 (.A1(\buffer[14][1][4] [13]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][4] [13]), .ZN(n_15_29_123));
   AOI22_X1 i_15_29_138 (.A1(\buffer[11][1][4] [13]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][4] [13]), .ZN(n_15_29_124));
   AOI22_X1 i_15_29_139 (.A1(\buffer[13][1][4] [13]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][1][4] [13]), .ZN(n_15_29_125));
   NAND4_X1 i_15_29_140 (.A1(n_15_29_134), .A2(n_15_29_132), .A3(n_15_29_130), 
      .A4(n_15_29_126), .ZN(\output_filter[1][4] [14]));
   AOI221_X1 i_15_29_141 (.A(n_15_29_127), .B1(n_25), .B2(\buffer[0][1][4] [14]), 
      .C1(\buffer[12][1][4] [14]), .C2(n_27), .ZN(n_15_29_126));
   NAND4_X1 i_15_29_142 (.A1(n_15_29_133), .A2(n_15_29_131), .A3(n_15_29_129), 
      .A4(n_15_29_128), .ZN(n_15_29_127));
   AOI22_X1 i_15_29_143 (.A1(\buffer[15][1][4] [14]), .A2(n_22), .B1(n_16), 
      .B2(\buffer[8][1][4] [14]), .ZN(n_15_29_128));
   AOI22_X1 i_15_29_144 (.A1(\buffer[10][1][4] [14]), .A2(n_21), .B1(n_29), 
      .B2(\buffer[7][1][4] [14]), .ZN(n_15_29_129));
   AOI22_X1 i_15_29_145 (.A1(\buffer[6][1][4] [14]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][4] [14]), .ZN(n_15_29_130));
   AOI22_X1 i_15_29_146 (.A1(\buffer[9][1][4] [14]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][4] [14]), .ZN(n_15_29_131));
   AOI22_X1 i_15_29_147 (.A1(\buffer[14][1][4] [14]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][4] [14]), .ZN(n_15_29_132));
   AOI22_X1 i_15_29_148 (.A1(\buffer[11][1][4] [14]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][4] [14]), .ZN(n_15_29_133));
   AOI22_X1 i_15_29_149 (.A1(\buffer[13][1][4] [14]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][4] [14]), .ZN(n_15_29_134));
   NAND2_X1 i_15_29_150 (.A1(n_15_29_137), .A2(n_15_29_135), .ZN(
      \output_filter[1][4] [15]));
   AOI221_X1 i_15_29_151 (.A(n_15_29_136), .B1(n_31), .B2(\buffer[3][1][4] [15]), 
      .C1(\buffer[14][1][4] [15]), .C2(n_19), .ZN(n_15_29_135));
   NAND3_X1 i_15_29_152 (.A1(n_15_29_143), .A2(n_15_29_141), .A3(n_15_29_139), 
      .ZN(n_15_29_136));
   AOI221_X1 i_15_29_153 (.A(n_15_29_138), .B1(n_16), .B2(\buffer[8][1][4] [15]), 
      .C1(\buffer[13][1][4] [15]), .C2(n_26), .ZN(n_15_29_137));
   NAND3_X1 i_15_29_154 (.A1(n_15_29_144), .A2(n_15_29_142), .A3(n_15_29_140), 
      .ZN(n_15_29_138));
   AOI22_X1 i_15_29_155 (.A1(\buffer[11][1][4] [15]), .A2(n_17), .B1(n_24), 
      .B2(\buffer[2][1][4] [15]), .ZN(n_15_29_139));
   AOI22_X1 i_15_29_156 (.A1(\buffer[10][1][4] [15]), .A2(n_21), .B1(n_23), 
      .B2(\buffer[1][1][4] [15]), .ZN(n_15_29_140));
   AOI22_X1 i_15_29_157 (.A1(\buffer[6][1][4] [15]), .A2(n_28), .B1(n_18), 
      .B2(\buffer[5][1][4] [15]), .ZN(n_15_29_141));
   AOI22_X1 i_15_29_158 (.A1(\buffer[9][1][4] [15]), .A2(n_20), .B1(n_30), 
      .B2(\buffer[4][1][4] [15]), .ZN(n_15_29_142));
   AOI22_X1 i_15_29_159 (.A1(\buffer[7][1][4] [15]), .A2(n_29), .B1(n_25), 
      .B2(\buffer[0][1][4] [15]), .ZN(n_15_29_143));
   AOI22_X1 i_15_29_160 (.A1(\buffer[15][1][4] [15]), .A2(n_22), .B1(n_27), 
      .B2(\buffer[12][1][4] [15]), .ZN(n_15_29_144));
   NAND4_X1 i_16_28_0 (.A1(n_16_28_8), .A2(n_16_28_6), .A3(n_16_28_4), .A4(
      n_16_28_0), .ZN(\output_filter[1][3] [0]));
   AOI221_X1 i_16_28_1 (.A(n_16_28_1), .B1(n_25), .B2(\buffer[0][1][3] [0]), 
      .C1(\buffer[12][1][3] [0]), .C2(n_27), .ZN(n_16_28_0));
   NAND4_X1 i_16_28_2 (.A1(n_16_28_7), .A2(n_16_28_5), .A3(n_16_28_3), .A4(
      n_16_28_2), .ZN(n_16_28_1));
   AOI22_X1 i_16_28_3 (.A1(\buffer[15][1][3] [0]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][3] [0]), .ZN(n_16_28_2));
   AOI22_X1 i_16_28_4 (.A1(\buffer[10][1][3] [0]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][3] [0]), .ZN(n_16_28_3));
   AOI22_X1 i_16_28_5 (.A1(\buffer[6][1][3] [0]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][1][3] [0]), .ZN(n_16_28_4));
   AOI22_X1 i_16_28_6 (.A1(\buffer[9][1][3] [0]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][1][3] [0]), .ZN(n_16_28_5));
   AOI22_X1 i_16_28_7 (.A1(\buffer[14][1][3] [0]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][3] [0]), .ZN(n_16_28_6));
   AOI22_X1 i_16_28_8 (.A1(\buffer[11][1][3] [0]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][3] [0]), .ZN(n_16_28_7));
   AOI22_X1 i_16_28_9 (.A1(\buffer[13][1][3] [0]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][3] [0]), .ZN(n_16_28_8));
   NAND4_X1 i_16_28_10 (.A1(n_16_28_17), .A2(n_16_28_15), .A3(n_16_28_13), 
      .A4(n_16_28_9), .ZN(\output_filter[1][3] [1]));
   AOI221_X1 i_16_28_11 (.A(n_16_28_10), .B1(n_25), .B2(\buffer[0][1][3] [1]), 
      .C1(\buffer[12][1][3] [1]), .C2(n_27), .ZN(n_16_28_9));
   NAND4_X1 i_16_28_12 (.A1(n_16_28_16), .A2(n_16_28_14), .A3(n_16_28_12), 
      .A4(n_16_28_11), .ZN(n_16_28_10));
   AOI22_X1 i_16_28_13 (.A1(\buffer[15][1][3] [1]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][3] [1]), .ZN(n_16_28_11));
   AOI22_X1 i_16_28_14 (.A1(\buffer[10][1][3] [1]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][3] [1]), .ZN(n_16_28_12));
   AOI22_X1 i_16_28_15 (.A1(\buffer[6][1][3] [1]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][3] [1]), .ZN(n_16_28_13));
   AOI22_X1 i_16_28_16 (.A1(\buffer[9][1][3] [1]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][3] [1]), .ZN(n_16_28_14));
   AOI22_X1 i_16_28_17 (.A1(\buffer[14][1][3] [1]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][3] [1]), .ZN(n_16_28_15));
   AOI22_X1 i_16_28_18 (.A1(\buffer[11][1][3] [1]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][3] [1]), .ZN(n_16_28_16));
   AOI22_X1 i_16_28_19 (.A1(\buffer[13][1][3] [1]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][3] [1]), .ZN(n_16_28_17));
   NAND4_X1 i_16_28_20 (.A1(n_16_28_26), .A2(n_16_28_24), .A3(n_16_28_22), 
      .A4(n_16_28_18), .ZN(\output_filter[1][3] [2]));
   AOI221_X1 i_16_28_21 (.A(n_16_28_19), .B1(n_25), .B2(\buffer[0][1][3] [2]), 
      .C1(\buffer[12][1][3] [2]), .C2(n_27), .ZN(n_16_28_18));
   NAND4_X1 i_16_28_22 (.A1(n_16_28_25), .A2(n_16_28_23), .A3(n_16_28_21), 
      .A4(n_16_28_20), .ZN(n_16_28_19));
   AOI22_X1 i_16_28_23 (.A1(\buffer[15][1][3] [2]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][3] [2]), .ZN(n_16_28_20));
   AOI22_X1 i_16_28_24 (.A1(\buffer[10][1][3] [2]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][3] [2]), .ZN(n_16_28_21));
   AOI22_X1 i_16_28_25 (.A1(\buffer[6][1][3] [2]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][3] [2]), .ZN(n_16_28_22));
   AOI22_X1 i_16_28_26 (.A1(\buffer[9][1][3] [2]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][3] [2]), .ZN(n_16_28_23));
   AOI22_X1 i_16_28_27 (.A1(\buffer[14][1][3] [2]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][3] [2]), .ZN(n_16_28_24));
   AOI22_X1 i_16_28_28 (.A1(\buffer[11][1][3] [2]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][3] [2]), .ZN(n_16_28_25));
   AOI22_X1 i_16_28_29 (.A1(\buffer[13][1][3] [2]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][3] [2]), .ZN(n_16_28_26));
   NAND4_X1 i_16_28_30 (.A1(n_16_28_35), .A2(n_16_28_33), .A3(n_16_28_31), 
      .A4(n_16_28_27), .ZN(\output_filter[1][3] [3]));
   AOI221_X1 i_16_28_31 (.A(n_16_28_28), .B1(n_25), .B2(\buffer[0][1][3] [3]), 
      .C1(\buffer[12][1][3] [3]), .C2(n_27), .ZN(n_16_28_27));
   NAND4_X1 i_16_28_32 (.A1(n_16_28_34), .A2(n_16_28_32), .A3(n_16_28_30), 
      .A4(n_16_28_29), .ZN(n_16_28_28));
   AOI22_X1 i_16_28_33 (.A1(\buffer[15][1][3] [3]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][3] [3]), .ZN(n_16_28_29));
   AOI22_X1 i_16_28_34 (.A1(\buffer[10][1][3] [3]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][3] [3]), .ZN(n_16_28_30));
   AOI22_X1 i_16_28_35 (.A1(\buffer[6][1][3] [3]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][3] [3]), .ZN(n_16_28_31));
   AOI22_X1 i_16_28_36 (.A1(\buffer[9][1][3] [3]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][3] [3]), .ZN(n_16_28_32));
   AOI22_X1 i_16_28_37 (.A1(\buffer[14][1][3] [3]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][3] [3]), .ZN(n_16_28_33));
   AOI22_X1 i_16_28_38 (.A1(\buffer[11][1][3] [3]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][3] [3]), .ZN(n_16_28_34));
   AOI22_X1 i_16_28_39 (.A1(\buffer[13][1][3] [3]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][3] [3]), .ZN(n_16_28_35));
   NAND4_X1 i_16_28_40 (.A1(n_16_28_44), .A2(n_16_28_42), .A3(n_16_28_40), 
      .A4(n_16_28_36), .ZN(\output_filter[1][3] [4]));
   AOI221_X1 i_16_28_41 (.A(n_16_28_37), .B1(n_25), .B2(\buffer[0][1][3] [4]), 
      .C1(\buffer[12][1][3] [4]), .C2(n_27), .ZN(n_16_28_36));
   NAND4_X1 i_16_28_42 (.A1(n_16_28_43), .A2(n_16_28_41), .A3(n_16_28_39), 
      .A4(n_16_28_38), .ZN(n_16_28_37));
   AOI22_X1 i_16_28_43 (.A1(\buffer[15][1][3] [4]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][3] [4]), .ZN(n_16_28_38));
   AOI22_X1 i_16_28_44 (.A1(\buffer[10][1][3] [4]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][3] [4]), .ZN(n_16_28_39));
   AOI22_X1 i_16_28_45 (.A1(\buffer[6][1][3] [4]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][3] [4]), .ZN(n_16_28_40));
   AOI22_X1 i_16_28_46 (.A1(\buffer[9][1][3] [4]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][1][3] [4]), .ZN(n_16_28_41));
   AOI22_X1 i_16_28_47 (.A1(\buffer[14][1][3] [4]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][3] [4]), .ZN(n_16_28_42));
   AOI22_X1 i_16_28_48 (.A1(\buffer[11][1][3] [4]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][3] [4]), .ZN(n_16_28_43));
   AOI22_X1 i_16_28_49 (.A1(\buffer[13][1][3] [4]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][1][3] [4]), .ZN(n_16_28_44));
   NAND4_X1 i_16_28_50 (.A1(n_16_28_53), .A2(n_16_28_51), .A3(n_16_28_49), 
      .A4(n_16_28_45), .ZN(\output_filter[1][3] [5]));
   AOI221_X1 i_16_28_51 (.A(n_16_28_46), .B1(n_25), .B2(\buffer[0][1][3] [5]), 
      .C1(\buffer[12][1][3] [5]), .C2(n_27), .ZN(n_16_28_45));
   NAND4_X1 i_16_28_52 (.A1(n_16_28_52), .A2(n_16_28_50), .A3(n_16_28_48), 
      .A4(n_16_28_47), .ZN(n_16_28_46));
   AOI22_X1 i_16_28_53 (.A1(\buffer[15][1][3] [5]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][3] [5]), .ZN(n_16_28_47));
   AOI22_X1 i_16_28_54 (.A1(\buffer[10][1][3] [5]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][3] [5]), .ZN(n_16_28_48));
   AOI22_X1 i_16_28_55 (.A1(\buffer[6][1][3] [5]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][3] [5]), .ZN(n_16_28_49));
   AOI22_X1 i_16_28_56 (.A1(\buffer[9][1][3] [5]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][3] [5]), .ZN(n_16_28_50));
   AOI22_X1 i_16_28_57 (.A1(\buffer[14][1][3] [5]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][3] [5]), .ZN(n_16_28_51));
   AOI22_X1 i_16_28_58 (.A1(\buffer[11][1][3] [5]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][3] [5]), .ZN(n_16_28_52));
   AOI22_X1 i_16_28_59 (.A1(\buffer[13][1][3] [5]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][3] [5]), .ZN(n_16_28_53));
   NAND4_X1 i_16_28_60 (.A1(n_16_28_62), .A2(n_16_28_60), .A3(n_16_28_58), 
      .A4(n_16_28_54), .ZN(\output_filter[1][3] [6]));
   AOI221_X1 i_16_28_61 (.A(n_16_28_55), .B1(n_25), .B2(\buffer[0][1][3] [6]), 
      .C1(\buffer[12][1][3] [6]), .C2(n_27), .ZN(n_16_28_54));
   NAND4_X1 i_16_28_62 (.A1(n_16_28_61), .A2(n_16_28_59), .A3(n_16_28_57), 
      .A4(n_16_28_56), .ZN(n_16_28_55));
   AOI22_X1 i_16_28_63 (.A1(\buffer[15][1][3] [6]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][3] [6]), .ZN(n_16_28_56));
   AOI22_X1 i_16_28_64 (.A1(\buffer[10][1][3] [6]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][3] [6]), .ZN(n_16_28_57));
   AOI22_X1 i_16_28_65 (.A1(\buffer[6][1][3] [6]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][3] [6]), .ZN(n_16_28_58));
   AOI22_X1 i_16_28_66 (.A1(\buffer[9][1][3] [6]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][3] [6]), .ZN(n_16_28_59));
   AOI22_X1 i_16_28_67 (.A1(\buffer[14][1][3] [6]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][3] [6]), .ZN(n_16_28_60));
   AOI22_X1 i_16_28_68 (.A1(\buffer[11][1][3] [6]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][3] [6]), .ZN(n_16_28_61));
   AOI22_X1 i_16_28_69 (.A1(\buffer[13][1][3] [6]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][3] [6]), .ZN(n_16_28_62));
   NAND4_X1 i_16_28_70 (.A1(n_16_28_71), .A2(n_16_28_69), .A3(n_16_28_67), 
      .A4(n_16_28_63), .ZN(\output_filter[1][3] [7]));
   AOI221_X1 i_16_28_71 (.A(n_16_28_64), .B1(n_25), .B2(\buffer[0][1][3] [7]), 
      .C1(\buffer[12][1][3] [7]), .C2(n_27), .ZN(n_16_28_63));
   NAND4_X1 i_16_28_72 (.A1(n_16_28_70), .A2(n_16_28_68), .A3(n_16_28_66), 
      .A4(n_16_28_65), .ZN(n_16_28_64));
   AOI22_X1 i_16_28_73 (.A1(\buffer[15][1][3] [7]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][3] [7]), .ZN(n_16_28_65));
   AOI22_X1 i_16_28_74 (.A1(\buffer[10][1][3] [7]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][3] [7]), .ZN(n_16_28_66));
   AOI22_X1 i_16_28_75 (.A1(\buffer[6][1][3] [7]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][3] [7]), .ZN(n_16_28_67));
   AOI22_X1 i_16_28_76 (.A1(\buffer[9][1][3] [7]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][1][3] [7]), .ZN(n_16_28_68));
   AOI22_X1 i_16_28_77 (.A1(\buffer[14][1][3] [7]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][3] [7]), .ZN(n_16_28_69));
   AOI22_X1 i_16_28_78 (.A1(\buffer[11][1][3] [7]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][3] [7]), .ZN(n_16_28_70));
   AOI22_X1 i_16_28_79 (.A1(\buffer[13][1][3] [7]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][1][3] [7]), .ZN(n_16_28_71));
   NAND4_X1 i_16_28_80 (.A1(n_16_28_80), .A2(n_16_28_78), .A3(n_16_28_76), 
      .A4(n_16_28_72), .ZN(\output_filter[1][3] [8]));
   AOI221_X1 i_16_28_81 (.A(n_16_28_73), .B1(n_25), .B2(\buffer[0][1][3] [8]), 
      .C1(\buffer[12][1][3] [8]), .C2(n_27), .ZN(n_16_28_72));
   NAND4_X1 i_16_28_82 (.A1(n_16_28_79), .A2(n_16_28_77), .A3(n_16_28_75), 
      .A4(n_16_28_74), .ZN(n_16_28_73));
   AOI22_X1 i_16_28_83 (.A1(\buffer[15][1][3] [8]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][3] [8]), .ZN(n_16_28_74));
   AOI22_X1 i_16_28_84 (.A1(\buffer[10][1][3] [8]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][3] [8]), .ZN(n_16_28_75));
   AOI22_X1 i_16_28_85 (.A1(\buffer[6][1][3] [8]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][3] [8]), .ZN(n_16_28_76));
   AOI22_X1 i_16_28_86 (.A1(\buffer[9][1][3] [8]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][3] [8]), .ZN(n_16_28_77));
   AOI22_X1 i_16_28_87 (.A1(\buffer[14][1][3] [8]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][3] [8]), .ZN(n_16_28_78));
   AOI22_X1 i_16_28_88 (.A1(\buffer[11][1][3] [8]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][3] [8]), .ZN(n_16_28_79));
   AOI22_X1 i_16_28_89 (.A1(\buffer[13][1][3] [8]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][3] [8]), .ZN(n_16_28_80));
   NAND4_X1 i_16_28_90 (.A1(n_16_28_89), .A2(n_16_28_87), .A3(n_16_28_85), 
      .A4(n_16_28_81), .ZN(\output_filter[1][3] [9]));
   AOI221_X1 i_16_28_91 (.A(n_16_28_82), .B1(n_25), .B2(\buffer[0][1][3] [9]), 
      .C1(\buffer[12][1][3] [9]), .C2(n_27), .ZN(n_16_28_81));
   NAND4_X1 i_16_28_92 (.A1(n_16_28_88), .A2(n_16_28_86), .A3(n_16_28_84), 
      .A4(n_16_28_83), .ZN(n_16_28_82));
   AOI22_X1 i_16_28_93 (.A1(\buffer[15][1][3] [9]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][3] [9]), .ZN(n_16_28_83));
   AOI22_X1 i_16_28_94 (.A1(\buffer[10][1][3] [9]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][3] [9]), .ZN(n_16_28_84));
   AOI22_X1 i_16_28_95 (.A1(\buffer[6][1][3] [9]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][3] [9]), .ZN(n_16_28_85));
   AOI22_X1 i_16_28_96 (.A1(\buffer[9][1][3] [9]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][1][3] [9]), .ZN(n_16_28_86));
   AOI22_X1 i_16_28_97 (.A1(\buffer[14][1][3] [9]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][3] [9]), .ZN(n_16_28_87));
   AOI22_X1 i_16_28_98 (.A1(\buffer[11][1][3] [9]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][3] [9]), .ZN(n_16_28_88));
   AOI22_X1 i_16_28_99 (.A1(\buffer[13][1][3] [9]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][1][3] [9]), .ZN(n_16_28_89));
   NAND4_X1 i_16_28_100 (.A1(n_16_28_98), .A2(n_16_28_96), .A3(n_16_28_94), 
      .A4(n_16_28_90), .ZN(\output_filter[1][3] [10]));
   AOI221_X1 i_16_28_101 (.A(n_16_28_91), .B1(n_25), .B2(\buffer[0][1][3] [10]), 
      .C1(\buffer[12][1][3] [10]), .C2(n_27), .ZN(n_16_28_90));
   NAND4_X1 i_16_28_102 (.A1(n_16_28_97), .A2(n_16_28_95), .A3(n_16_28_93), 
      .A4(n_16_28_92), .ZN(n_16_28_91));
   AOI22_X1 i_16_28_103 (.A1(\buffer[15][1][3] [10]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][3] [10]), .ZN(n_16_28_92));
   AOI22_X1 i_16_28_104 (.A1(\buffer[10][1][3] [10]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][3] [10]), .ZN(n_16_28_93));
   AOI22_X1 i_16_28_105 (.A1(\buffer[6][1][3] [10]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][3] [10]), .ZN(n_16_28_94));
   AOI22_X1 i_16_28_106 (.A1(\buffer[9][1][3] [10]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][3] [10]), .ZN(n_16_28_95));
   AOI22_X1 i_16_28_107 (.A1(\buffer[14][1][3] [10]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][3] [10]), .ZN(n_16_28_96));
   AOI22_X1 i_16_28_108 (.A1(\buffer[11][1][3] [10]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][3] [10]), .ZN(n_16_28_97));
   AOI22_X1 i_16_28_109 (.A1(\buffer[13][1][3] [10]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][3] [10]), .ZN(n_16_28_98));
   NAND4_X1 i_16_28_110 (.A1(n_16_28_107), .A2(n_16_28_105), .A3(n_16_28_103), 
      .A4(n_16_28_99), .ZN(\output_filter[1][3] [11]));
   AOI221_X1 i_16_28_111 (.A(n_16_28_100), .B1(n_25), .B2(\buffer[0][1][3] [11]), 
      .C1(\buffer[12][1][3] [11]), .C2(n_27), .ZN(n_16_28_99));
   NAND4_X1 i_16_28_112 (.A1(n_16_28_106), .A2(n_16_28_104), .A3(n_16_28_102), 
      .A4(n_16_28_101), .ZN(n_16_28_100));
   AOI22_X1 i_16_28_113 (.A1(\buffer[15][1][3] [11]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][3] [11]), .ZN(n_16_28_101));
   AOI22_X1 i_16_28_114 (.A1(\buffer[10][1][3] [11]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][3] [11]), .ZN(n_16_28_102));
   AOI22_X1 i_16_28_115 (.A1(\buffer[6][1][3] [11]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][3] [11]), .ZN(n_16_28_103));
   AOI22_X1 i_16_28_116 (.A1(\buffer[9][1][3] [11]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][1][3] [11]), .ZN(n_16_28_104));
   AOI22_X1 i_16_28_117 (.A1(\buffer[14][1][3] [11]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][3] [11]), .ZN(n_16_28_105));
   AOI22_X1 i_16_28_118 (.A1(\buffer[11][1][3] [11]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][3] [11]), .ZN(n_16_28_106));
   AOI22_X1 i_16_28_119 (.A1(\buffer[13][1][3] [11]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][1][3] [11]), .ZN(n_16_28_107));
   NAND4_X1 i_16_28_120 (.A1(n_16_28_116), .A2(n_16_28_114), .A3(n_16_28_112), 
      .A4(n_16_28_108), .ZN(\output_filter[1][3] [12]));
   AOI221_X1 i_16_28_121 (.A(n_16_28_109), .B1(n_25), .B2(\buffer[0][1][3] [12]), 
      .C1(\buffer[12][1][3] [12]), .C2(n_27), .ZN(n_16_28_108));
   NAND4_X1 i_16_28_122 (.A1(n_16_28_115), .A2(n_16_28_113), .A3(n_16_28_111), 
      .A4(n_16_28_110), .ZN(n_16_28_109));
   AOI22_X1 i_16_28_123 (.A1(\buffer[15][1][3] [12]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][3] [12]), .ZN(n_16_28_110));
   AOI22_X1 i_16_28_124 (.A1(\buffer[10][1][3] [12]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][3] [12]), .ZN(n_16_28_111));
   AOI22_X1 i_16_28_125 (.A1(\buffer[6][1][3] [12]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][3] [12]), .ZN(n_16_28_112));
   AOI22_X1 i_16_28_126 (.A1(\buffer[9][1][3] [12]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][3] [12]), .ZN(n_16_28_113));
   AOI22_X1 i_16_28_127 (.A1(\buffer[14][1][3] [12]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][3] [12]), .ZN(n_16_28_114));
   AOI22_X1 i_16_28_128 (.A1(\buffer[11][1][3] [12]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][3] [12]), .ZN(n_16_28_115));
   AOI22_X1 i_16_28_129 (.A1(\buffer[13][1][3] [12]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][3] [12]), .ZN(n_16_28_116));
   NAND4_X1 i_16_28_130 (.A1(n_16_28_125), .A2(n_16_28_123), .A3(n_16_28_121), 
      .A4(n_16_28_117), .ZN(\output_filter[1][3] [13]));
   AOI221_X1 i_16_28_131 (.A(n_16_28_118), .B1(n_25), .B2(\buffer[0][1][3] [13]), 
      .C1(\buffer[12][1][3] [13]), .C2(n_27), .ZN(n_16_28_117));
   NAND4_X1 i_16_28_132 (.A1(n_16_28_124), .A2(n_16_28_122), .A3(n_16_28_120), 
      .A4(n_16_28_119), .ZN(n_16_28_118));
   AOI22_X1 i_16_28_133 (.A1(\buffer[15][1][3] [13]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][3] [13]), .ZN(n_16_28_119));
   AOI22_X1 i_16_28_134 (.A1(\buffer[10][1][3] [13]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][3] [13]), .ZN(n_16_28_120));
   AOI22_X1 i_16_28_135 (.A1(\buffer[6][1][3] [13]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][3] [13]), .ZN(n_16_28_121));
   AOI22_X1 i_16_28_136 (.A1(\buffer[9][1][3] [13]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][1][3] [13]), .ZN(n_16_28_122));
   AOI22_X1 i_16_28_137 (.A1(\buffer[14][1][3] [13]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][3] [13]), .ZN(n_16_28_123));
   AOI22_X1 i_16_28_138 (.A1(\buffer[11][1][3] [13]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][3] [13]), .ZN(n_16_28_124));
   AOI22_X1 i_16_28_139 (.A1(\buffer[13][1][3] [13]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][1][3] [13]), .ZN(n_16_28_125));
   NAND4_X1 i_16_28_140 (.A1(n_16_28_134), .A2(n_16_28_132), .A3(n_16_28_130), 
      .A4(n_16_28_126), .ZN(\output_filter[1][3] [14]));
   AOI221_X1 i_16_28_141 (.A(n_16_28_127), .B1(n_25), .B2(\buffer[0][1][3] [14]), 
      .C1(\buffer[12][1][3] [14]), .C2(n_27), .ZN(n_16_28_126));
   NAND4_X1 i_16_28_142 (.A1(n_16_28_133), .A2(n_16_28_131), .A3(n_16_28_129), 
      .A4(n_16_28_128), .ZN(n_16_28_127));
   AOI22_X1 i_16_28_143 (.A1(\buffer[15][1][3] [14]), .A2(n_22), .B1(n_16), 
      .B2(\buffer[8][1][3] [14]), .ZN(n_16_28_128));
   AOI22_X1 i_16_28_144 (.A1(\buffer[10][1][3] [14]), .A2(n_21), .B1(n_29), 
      .B2(\buffer[7][1][3] [14]), .ZN(n_16_28_129));
   AOI22_X1 i_16_28_145 (.A1(\buffer[6][1][3] [14]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][3] [14]), .ZN(n_16_28_130));
   AOI22_X1 i_16_28_146 (.A1(\buffer[9][1][3] [14]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][3] [14]), .ZN(n_16_28_131));
   AOI22_X1 i_16_28_147 (.A1(\buffer[14][1][3] [14]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][3] [14]), .ZN(n_16_28_132));
   AOI22_X1 i_16_28_148 (.A1(\buffer[11][1][3] [14]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][3] [14]), .ZN(n_16_28_133));
   AOI22_X1 i_16_28_149 (.A1(\buffer[13][1][3] [14]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][3] [14]), .ZN(n_16_28_134));
   NAND2_X1 i_16_28_150 (.A1(n_16_28_137), .A2(n_16_28_135), .ZN(
      \output_filter[1][3] [15]));
   AOI221_X1 i_16_28_151 (.A(n_16_28_136), .B1(n_31), .B2(\buffer[3][1][3] [15]), 
      .C1(\buffer[14][1][3] [15]), .C2(n_19), .ZN(n_16_28_135));
   NAND3_X1 i_16_28_152 (.A1(n_16_28_143), .A2(n_16_28_141), .A3(n_16_28_139), 
      .ZN(n_16_28_136));
   AOI221_X1 i_16_28_153 (.A(n_16_28_138), .B1(n_16), .B2(\buffer[8][1][3] [15]), 
      .C1(\buffer[13][1][3] [15]), .C2(n_26), .ZN(n_16_28_137));
   NAND3_X1 i_16_28_154 (.A1(n_16_28_144), .A2(n_16_28_142), .A3(n_16_28_140), 
      .ZN(n_16_28_138));
   AOI22_X1 i_16_28_155 (.A1(\buffer[11][1][3] [15]), .A2(n_17), .B1(n_24), 
      .B2(\buffer[2][1][3] [15]), .ZN(n_16_28_139));
   AOI22_X1 i_16_28_156 (.A1(\buffer[10][1][3] [15]), .A2(n_21), .B1(n_23), 
      .B2(\buffer[1][1][3] [15]), .ZN(n_16_28_140));
   AOI22_X1 i_16_28_157 (.A1(\buffer[6][1][3] [15]), .A2(n_28), .B1(n_18), 
      .B2(\buffer[5][1][3] [15]), .ZN(n_16_28_141));
   AOI22_X1 i_16_28_158 (.A1(\buffer[9][1][3] [15]), .A2(n_20), .B1(n_30), 
      .B2(\buffer[4][1][3] [15]), .ZN(n_16_28_142));
   AOI22_X1 i_16_28_159 (.A1(\buffer[7][1][3] [15]), .A2(n_29), .B1(n_25), 
      .B2(\buffer[0][1][3] [15]), .ZN(n_16_28_143));
   AOI22_X1 i_16_28_160 (.A1(\buffer[15][1][3] [15]), .A2(n_22), .B1(n_27), 
      .B2(\buffer[12][1][3] [15]), .ZN(n_16_28_144));
   NAND4_X1 i_17_34_0 (.A1(n_17_34_8), .A2(n_17_34_6), .A3(n_17_34_4), .A4(
      n_17_34_0), .ZN(\output_filter[2][4] [0]));
   AOI221_X1 i_17_34_1 (.A(n_17_34_1), .B1(n_25), .B2(\buffer[0][2][4] [0]), 
      .C1(\buffer[12][2][4] [0]), .C2(n_27), .ZN(n_17_34_0));
   NAND4_X1 i_17_34_2 (.A1(n_17_34_7), .A2(n_17_34_5), .A3(n_17_34_3), .A4(
      n_17_34_2), .ZN(n_17_34_1));
   AOI22_X1 i_17_34_3 (.A1(\buffer[15][2][4] [0]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][4] [0]), .ZN(n_17_34_2));
   AOI22_X1 i_17_34_4 (.A1(\buffer[10][2][4] [0]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][4] [0]), .ZN(n_17_34_3));
   AOI22_X1 i_17_34_5 (.A1(\buffer[6][2][4] [0]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][2][4] [0]), .ZN(n_17_34_4));
   AOI22_X1 i_17_34_6 (.A1(\buffer[9][2][4] [0]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][2][4] [0]), .ZN(n_17_34_5));
   AOI22_X1 i_17_34_7 (.A1(\buffer[14][2][4] [0]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][4] [0]), .ZN(n_17_34_6));
   AOI22_X1 i_17_34_8 (.A1(\buffer[11][2][4] [0]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][4] [0]), .ZN(n_17_34_7));
   AOI22_X1 i_17_34_9 (.A1(\buffer[13][2][4] [0]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][4] [0]), .ZN(n_17_34_8));
   NAND4_X1 i_17_34_10 (.A1(n_17_34_17), .A2(n_17_34_15), .A3(n_17_34_13), 
      .A4(n_17_34_9), .ZN(\output_filter[2][4] [1]));
   AOI221_X1 i_17_34_11 (.A(n_17_34_10), .B1(n_25), .B2(\buffer[0][2][4] [1]), 
      .C1(\buffer[12][2][4] [1]), .C2(n_27), .ZN(n_17_34_9));
   NAND4_X1 i_17_34_12 (.A1(n_17_34_16), .A2(n_17_34_14), .A3(n_17_34_12), 
      .A4(n_17_34_11), .ZN(n_17_34_10));
   AOI22_X1 i_17_34_13 (.A1(\buffer[15][2][4] [1]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][4] [1]), .ZN(n_17_34_11));
   AOI22_X1 i_17_34_14 (.A1(\buffer[10][2][4] [1]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][4] [1]), .ZN(n_17_34_12));
   AOI22_X1 i_17_34_15 (.A1(\buffer[6][2][4] [1]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][4] [1]), .ZN(n_17_34_13));
   AOI22_X1 i_17_34_16 (.A1(\buffer[9][2][4] [1]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][4] [1]), .ZN(n_17_34_14));
   AOI22_X1 i_17_34_17 (.A1(\buffer[14][2][4] [1]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][4] [1]), .ZN(n_17_34_15));
   AOI22_X1 i_17_34_18 (.A1(\buffer[11][2][4] [1]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][4] [1]), .ZN(n_17_34_16));
   AOI22_X1 i_17_34_19 (.A1(\buffer[13][2][4] [1]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][4] [1]), .ZN(n_17_34_17));
   NAND4_X1 i_17_34_20 (.A1(n_17_34_26), .A2(n_17_34_24), .A3(n_17_34_22), 
      .A4(n_17_34_18), .ZN(\output_filter[2][4] [2]));
   AOI221_X1 i_17_34_21 (.A(n_17_34_19), .B1(n_25), .B2(\buffer[0][2][4] [2]), 
      .C1(\buffer[12][2][4] [2]), .C2(n_27), .ZN(n_17_34_18));
   NAND4_X1 i_17_34_22 (.A1(n_17_34_25), .A2(n_17_34_23), .A3(n_17_34_21), 
      .A4(n_17_34_20), .ZN(n_17_34_19));
   AOI22_X1 i_17_34_23 (.A1(\buffer[15][2][4] [2]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][4] [2]), .ZN(n_17_34_20));
   AOI22_X1 i_17_34_24 (.A1(\buffer[10][2][4] [2]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][4] [2]), .ZN(n_17_34_21));
   AOI22_X1 i_17_34_25 (.A1(\buffer[6][2][4] [2]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][4] [2]), .ZN(n_17_34_22));
   AOI22_X1 i_17_34_26 (.A1(\buffer[9][2][4] [2]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][4] [2]), .ZN(n_17_34_23));
   AOI22_X1 i_17_34_27 (.A1(\buffer[14][2][4] [2]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][4] [2]), .ZN(n_17_34_24));
   AOI22_X1 i_17_34_28 (.A1(\buffer[11][2][4] [2]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][4] [2]), .ZN(n_17_34_25));
   AOI22_X1 i_17_34_29 (.A1(\buffer[13][2][4] [2]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][4] [2]), .ZN(n_17_34_26));
   NAND4_X1 i_17_34_30 (.A1(n_17_34_35), .A2(n_17_34_33), .A3(n_17_34_31), 
      .A4(n_17_34_27), .ZN(\output_filter[2][4] [3]));
   AOI221_X1 i_17_34_31 (.A(n_17_34_28), .B1(n_25), .B2(\buffer[0][2][4] [3]), 
      .C1(\buffer[12][2][4] [3]), .C2(n_27), .ZN(n_17_34_27));
   NAND4_X1 i_17_34_32 (.A1(n_17_34_34), .A2(n_17_34_32), .A3(n_17_34_30), 
      .A4(n_17_34_29), .ZN(n_17_34_28));
   AOI22_X1 i_17_34_33 (.A1(\buffer[15][2][4] [3]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][4] [3]), .ZN(n_17_34_29));
   AOI22_X1 i_17_34_34 (.A1(\buffer[10][2][4] [3]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][4] [3]), .ZN(n_17_34_30));
   AOI22_X1 i_17_34_35 (.A1(\buffer[6][2][4] [3]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][4] [3]), .ZN(n_17_34_31));
   AOI22_X1 i_17_34_36 (.A1(\buffer[9][2][4] [3]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][4] [3]), .ZN(n_17_34_32));
   AOI22_X1 i_17_34_37 (.A1(\buffer[14][2][4] [3]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][4] [3]), .ZN(n_17_34_33));
   AOI22_X1 i_17_34_38 (.A1(\buffer[11][2][4] [3]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][4] [3]), .ZN(n_17_34_34));
   AOI22_X1 i_17_34_39 (.A1(\buffer[13][2][4] [3]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][4] [3]), .ZN(n_17_34_35));
   NAND4_X1 i_17_34_40 (.A1(n_17_34_44), .A2(n_17_34_42), .A3(n_17_34_40), 
      .A4(n_17_34_36), .ZN(\output_filter[2][4] [4]));
   AOI221_X1 i_17_34_41 (.A(n_17_34_37), .B1(n_25), .B2(\buffer[0][2][4] [4]), 
      .C1(\buffer[12][2][4] [4]), .C2(n_27), .ZN(n_17_34_36));
   NAND4_X1 i_17_34_42 (.A1(n_17_34_43), .A2(n_17_34_41), .A3(n_17_34_39), 
      .A4(n_17_34_38), .ZN(n_17_34_37));
   AOI22_X1 i_17_34_43 (.A1(\buffer[15][2][4] [4]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][4] [4]), .ZN(n_17_34_38));
   AOI22_X1 i_17_34_44 (.A1(\buffer[10][2][4] [4]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][4] [4]), .ZN(n_17_34_39));
   AOI22_X1 i_17_34_45 (.A1(\buffer[6][2][4] [4]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][4] [4]), .ZN(n_17_34_40));
   AOI22_X1 i_17_34_46 (.A1(\buffer[9][2][4] [4]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][2][4] [4]), .ZN(n_17_34_41));
   AOI22_X1 i_17_34_47 (.A1(\buffer[14][2][4] [4]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][4] [4]), .ZN(n_17_34_42));
   AOI22_X1 i_17_34_48 (.A1(\buffer[11][2][4] [4]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][4] [4]), .ZN(n_17_34_43));
   AOI22_X1 i_17_34_49 (.A1(\buffer[13][2][4] [4]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][2][4] [4]), .ZN(n_17_34_44));
   NAND4_X1 i_17_34_50 (.A1(n_17_34_53), .A2(n_17_34_51), .A3(n_17_34_49), 
      .A4(n_17_34_45), .ZN(\output_filter[2][4] [5]));
   AOI221_X1 i_17_34_51 (.A(n_17_34_46), .B1(n_25), .B2(\buffer[0][2][4] [5]), 
      .C1(\buffer[12][2][4] [5]), .C2(n_27), .ZN(n_17_34_45));
   NAND4_X1 i_17_34_52 (.A1(n_17_34_52), .A2(n_17_34_50), .A3(n_17_34_48), 
      .A4(n_17_34_47), .ZN(n_17_34_46));
   AOI22_X1 i_17_34_53 (.A1(\buffer[15][2][4] [5]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][4] [5]), .ZN(n_17_34_47));
   AOI22_X1 i_17_34_54 (.A1(\buffer[10][2][4] [5]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][4] [5]), .ZN(n_17_34_48));
   AOI22_X1 i_17_34_55 (.A1(\buffer[6][2][4] [5]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][4] [5]), .ZN(n_17_34_49));
   AOI22_X1 i_17_34_56 (.A1(\buffer[9][2][4] [5]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][4] [5]), .ZN(n_17_34_50));
   AOI22_X1 i_17_34_57 (.A1(\buffer[14][2][4] [5]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][4] [5]), .ZN(n_17_34_51));
   AOI22_X1 i_17_34_58 (.A1(\buffer[11][2][4] [5]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][4] [5]), .ZN(n_17_34_52));
   AOI22_X1 i_17_34_59 (.A1(\buffer[13][2][4] [5]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][4] [5]), .ZN(n_17_34_53));
   NAND4_X1 i_17_34_60 (.A1(n_17_34_62), .A2(n_17_34_60), .A3(n_17_34_58), 
      .A4(n_17_34_54), .ZN(\output_filter[2][4] [6]));
   AOI221_X1 i_17_34_61 (.A(n_17_34_55), .B1(n_25), .B2(\buffer[0][2][4] [6]), 
      .C1(\buffer[12][2][4] [6]), .C2(n_27), .ZN(n_17_34_54));
   NAND4_X1 i_17_34_62 (.A1(n_17_34_61), .A2(n_17_34_59), .A3(n_17_34_57), 
      .A4(n_17_34_56), .ZN(n_17_34_55));
   AOI22_X1 i_17_34_63 (.A1(\buffer[15][2][4] [6]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][4] [6]), .ZN(n_17_34_56));
   AOI22_X1 i_17_34_64 (.A1(\buffer[10][2][4] [6]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][4] [6]), .ZN(n_17_34_57));
   AOI22_X1 i_17_34_65 (.A1(\buffer[6][2][4] [6]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][4] [6]), .ZN(n_17_34_58));
   AOI22_X1 i_17_34_66 (.A1(\buffer[9][2][4] [6]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][4] [6]), .ZN(n_17_34_59));
   AOI22_X1 i_17_34_67 (.A1(\buffer[14][2][4] [6]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][4] [6]), .ZN(n_17_34_60));
   AOI22_X1 i_17_34_68 (.A1(\buffer[11][2][4] [6]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][4] [6]), .ZN(n_17_34_61));
   AOI22_X1 i_17_34_69 (.A1(\buffer[13][2][4] [6]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][4] [6]), .ZN(n_17_34_62));
   NAND4_X1 i_17_34_70 (.A1(n_17_34_71), .A2(n_17_34_69), .A3(n_17_34_67), 
      .A4(n_17_34_63), .ZN(\output_filter[2][4] [7]));
   AOI221_X1 i_17_34_71 (.A(n_17_34_64), .B1(n_25), .B2(\buffer[0][2][4] [7]), 
      .C1(\buffer[12][2][4] [7]), .C2(n_27), .ZN(n_17_34_63));
   NAND4_X1 i_17_34_72 (.A1(n_17_34_70), .A2(n_17_34_68), .A3(n_17_34_66), 
      .A4(n_17_34_65), .ZN(n_17_34_64));
   AOI22_X1 i_17_34_73 (.A1(\buffer[15][2][4] [7]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][4] [7]), .ZN(n_17_34_65));
   AOI22_X1 i_17_34_74 (.A1(\buffer[10][2][4] [7]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][4] [7]), .ZN(n_17_34_66));
   AOI22_X1 i_17_34_75 (.A1(\buffer[6][2][4] [7]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][4] [7]), .ZN(n_17_34_67));
   AOI22_X1 i_17_34_76 (.A1(\buffer[9][2][4] [7]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][2][4] [7]), .ZN(n_17_34_68));
   AOI22_X1 i_17_34_77 (.A1(\buffer[14][2][4] [7]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][4] [7]), .ZN(n_17_34_69));
   AOI22_X1 i_17_34_78 (.A1(\buffer[11][2][4] [7]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][4] [7]), .ZN(n_17_34_70));
   AOI22_X1 i_17_34_79 (.A1(\buffer[13][2][4] [7]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][2][4] [7]), .ZN(n_17_34_71));
   NAND4_X1 i_17_34_80 (.A1(n_17_34_80), .A2(n_17_34_78), .A3(n_17_34_76), 
      .A4(n_17_34_72), .ZN(\output_filter[2][4] [8]));
   AOI221_X1 i_17_34_81 (.A(n_17_34_73), .B1(n_25), .B2(\buffer[0][2][4] [8]), 
      .C1(\buffer[12][2][4] [8]), .C2(n_27), .ZN(n_17_34_72));
   NAND4_X1 i_17_34_82 (.A1(n_17_34_79), .A2(n_17_34_77), .A3(n_17_34_75), 
      .A4(n_17_34_74), .ZN(n_17_34_73));
   AOI22_X1 i_17_34_83 (.A1(\buffer[15][2][4] [8]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][4] [8]), .ZN(n_17_34_74));
   AOI22_X1 i_17_34_84 (.A1(\buffer[10][2][4] [8]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][4] [8]), .ZN(n_17_34_75));
   AOI22_X1 i_17_34_85 (.A1(\buffer[6][2][4] [8]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][4] [8]), .ZN(n_17_34_76));
   AOI22_X1 i_17_34_86 (.A1(\buffer[9][2][4] [8]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][4] [8]), .ZN(n_17_34_77));
   AOI22_X1 i_17_34_87 (.A1(\buffer[14][2][4] [8]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][4] [8]), .ZN(n_17_34_78));
   AOI22_X1 i_17_34_88 (.A1(\buffer[11][2][4] [8]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][4] [8]), .ZN(n_17_34_79));
   AOI22_X1 i_17_34_89 (.A1(\buffer[13][2][4] [8]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][4] [8]), .ZN(n_17_34_80));
   NAND4_X1 i_17_34_90 (.A1(n_17_34_89), .A2(n_17_34_87), .A3(n_17_34_85), 
      .A4(n_17_34_81), .ZN(\output_filter[2][4] [9]));
   AOI221_X1 i_17_34_91 (.A(n_17_34_82), .B1(n_25), .B2(\buffer[0][2][4] [9]), 
      .C1(\buffer[12][2][4] [9]), .C2(n_27), .ZN(n_17_34_81));
   NAND4_X1 i_17_34_92 (.A1(n_17_34_88), .A2(n_17_34_86), .A3(n_17_34_84), 
      .A4(n_17_34_83), .ZN(n_17_34_82));
   AOI22_X1 i_17_34_93 (.A1(\buffer[15][2][4] [9]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][4] [9]), .ZN(n_17_34_83));
   AOI22_X1 i_17_34_94 (.A1(\buffer[10][2][4] [9]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][4] [9]), .ZN(n_17_34_84));
   AOI22_X1 i_17_34_95 (.A1(\buffer[6][2][4] [9]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][4] [9]), .ZN(n_17_34_85));
   AOI22_X1 i_17_34_96 (.A1(\buffer[9][2][4] [9]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][2][4] [9]), .ZN(n_17_34_86));
   AOI22_X1 i_17_34_97 (.A1(\buffer[14][2][4] [9]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][4] [9]), .ZN(n_17_34_87));
   AOI22_X1 i_17_34_98 (.A1(\buffer[11][2][4] [9]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][4] [9]), .ZN(n_17_34_88));
   AOI22_X1 i_17_34_99 (.A1(\buffer[13][2][4] [9]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][2][4] [9]), .ZN(n_17_34_89));
   NAND4_X1 i_17_34_100 (.A1(n_17_34_98), .A2(n_17_34_96), .A3(n_17_34_94), 
      .A4(n_17_34_90), .ZN(\output_filter[2][4] [10]));
   AOI221_X1 i_17_34_101 (.A(n_17_34_91), .B1(n_25), .B2(\buffer[0][2][4] [10]), 
      .C1(\buffer[12][2][4] [10]), .C2(n_27), .ZN(n_17_34_90));
   NAND4_X1 i_17_34_102 (.A1(n_17_34_97), .A2(n_17_34_95), .A3(n_17_34_93), 
      .A4(n_17_34_92), .ZN(n_17_34_91));
   AOI22_X1 i_17_34_103 (.A1(\buffer[15][2][4] [10]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][4] [10]), .ZN(n_17_34_92));
   AOI22_X1 i_17_34_104 (.A1(\buffer[10][2][4] [10]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][4] [10]), .ZN(n_17_34_93));
   AOI22_X1 i_17_34_105 (.A1(\buffer[6][2][4] [10]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][4] [10]), .ZN(n_17_34_94));
   AOI22_X1 i_17_34_106 (.A1(\buffer[9][2][4] [10]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][4] [10]), .ZN(n_17_34_95));
   AOI22_X1 i_17_34_107 (.A1(\buffer[14][2][4] [10]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][4] [10]), .ZN(n_17_34_96));
   AOI22_X1 i_17_34_108 (.A1(\buffer[11][2][4] [10]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][4] [10]), .ZN(n_17_34_97));
   AOI22_X1 i_17_34_109 (.A1(\buffer[13][2][4] [10]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][4] [10]), .ZN(n_17_34_98));
   NAND4_X1 i_17_34_110 (.A1(n_17_34_107), .A2(n_17_34_105), .A3(n_17_34_103), 
      .A4(n_17_34_99), .ZN(\output_filter[2][4] [11]));
   AOI221_X1 i_17_34_111 (.A(n_17_34_100), .B1(n_25), .B2(\buffer[0][2][4] [11]), 
      .C1(\buffer[12][2][4] [11]), .C2(n_27), .ZN(n_17_34_99));
   NAND4_X1 i_17_34_112 (.A1(n_17_34_106), .A2(n_17_34_104), .A3(n_17_34_102), 
      .A4(n_17_34_101), .ZN(n_17_34_100));
   AOI22_X1 i_17_34_113 (.A1(\buffer[15][2][4] [11]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][4] [11]), .ZN(n_17_34_101));
   AOI22_X1 i_17_34_114 (.A1(\buffer[10][2][4] [11]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][4] [11]), .ZN(n_17_34_102));
   AOI22_X1 i_17_34_115 (.A1(\buffer[6][2][4] [11]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][4] [11]), .ZN(n_17_34_103));
   AOI22_X1 i_17_34_116 (.A1(\buffer[9][2][4] [11]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][2][4] [11]), .ZN(n_17_34_104));
   AOI22_X1 i_17_34_117 (.A1(\buffer[14][2][4] [11]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][4] [11]), .ZN(n_17_34_105));
   AOI22_X1 i_17_34_118 (.A1(\buffer[11][2][4] [11]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][4] [11]), .ZN(n_17_34_106));
   AOI22_X1 i_17_34_119 (.A1(\buffer[13][2][4] [11]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][2][4] [11]), .ZN(n_17_34_107));
   NAND4_X1 i_17_34_120 (.A1(n_17_34_116), .A2(n_17_34_114), .A3(n_17_34_112), 
      .A4(n_17_34_108), .ZN(\output_filter[2][4] [12]));
   AOI221_X1 i_17_34_121 (.A(n_17_34_109), .B1(n_25), .B2(\buffer[0][2][4] [12]), 
      .C1(\buffer[12][2][4] [12]), .C2(n_27), .ZN(n_17_34_108));
   NAND4_X1 i_17_34_122 (.A1(n_17_34_115), .A2(n_17_34_113), .A3(n_17_34_111), 
      .A4(n_17_34_110), .ZN(n_17_34_109));
   AOI22_X1 i_17_34_123 (.A1(\buffer[15][2][4] [12]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][4] [12]), .ZN(n_17_34_110));
   AOI22_X1 i_17_34_124 (.A1(\buffer[10][2][4] [12]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][4] [12]), .ZN(n_17_34_111));
   AOI22_X1 i_17_34_125 (.A1(\buffer[6][2][4] [12]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][4] [12]), .ZN(n_17_34_112));
   AOI22_X1 i_17_34_126 (.A1(\buffer[9][2][4] [12]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][4] [12]), .ZN(n_17_34_113));
   AOI22_X1 i_17_34_127 (.A1(\buffer[14][2][4] [12]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][4] [12]), .ZN(n_17_34_114));
   AOI22_X1 i_17_34_128 (.A1(\buffer[11][2][4] [12]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][4] [12]), .ZN(n_17_34_115));
   AOI22_X1 i_17_34_129 (.A1(\buffer[13][2][4] [12]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][4] [12]), .ZN(n_17_34_116));
   NAND4_X1 i_17_34_130 (.A1(n_17_34_125), .A2(n_17_34_123), .A3(n_17_34_121), 
      .A4(n_17_34_117), .ZN(\output_filter[2][4] [13]));
   AOI221_X1 i_17_34_131 (.A(n_17_34_118), .B1(n_25), .B2(\buffer[0][2][4] [13]), 
      .C1(\buffer[12][2][4] [13]), .C2(n_27), .ZN(n_17_34_117));
   NAND4_X1 i_17_34_132 (.A1(n_17_34_124), .A2(n_17_34_122), .A3(n_17_34_120), 
      .A4(n_17_34_119), .ZN(n_17_34_118));
   AOI22_X1 i_17_34_133 (.A1(\buffer[15][2][4] [13]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][2][4] [13]), .ZN(n_17_34_119));
   AOI22_X1 i_17_34_134 (.A1(\buffer[10][2][4] [13]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][2][4] [13]), .ZN(n_17_34_120));
   AOI22_X1 i_17_34_135 (.A1(\buffer[6][2][4] [13]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][4] [13]), .ZN(n_17_34_121));
   AOI22_X1 i_17_34_136 (.A1(\buffer[9][2][4] [13]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][2][4] [13]), .ZN(n_17_34_122));
   AOI22_X1 i_17_34_137 (.A1(\buffer[14][2][4] [13]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][4] [13]), .ZN(n_17_34_123));
   AOI22_X1 i_17_34_138 (.A1(\buffer[11][2][4] [13]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][4] [13]), .ZN(n_17_34_124));
   AOI22_X1 i_17_34_139 (.A1(\buffer[13][2][4] [13]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][2][4] [13]), .ZN(n_17_34_125));
   NAND4_X1 i_17_34_140 (.A1(n_17_34_134), .A2(n_17_34_132), .A3(n_17_34_130), 
      .A4(n_17_34_126), .ZN(\output_filter[2][4] [14]));
   AOI221_X1 i_17_34_141 (.A(n_17_34_127), .B1(n_25), .B2(\buffer[0][2][4] [14]), 
      .C1(\buffer[12][2][4] [14]), .C2(n_27), .ZN(n_17_34_126));
   NAND4_X1 i_17_34_142 (.A1(n_17_34_133), .A2(n_17_34_131), .A3(n_17_34_129), 
      .A4(n_17_34_128), .ZN(n_17_34_127));
   AOI22_X1 i_17_34_143 (.A1(\buffer[15][2][4] [14]), .A2(n_22), .B1(n_16), 
      .B2(\buffer[8][2][4] [14]), .ZN(n_17_34_128));
   AOI22_X1 i_17_34_144 (.A1(\buffer[10][2][4] [14]), .A2(n_21), .B1(n_29), 
      .B2(\buffer[7][2][4] [14]), .ZN(n_17_34_129));
   AOI22_X1 i_17_34_145 (.A1(\buffer[6][2][4] [14]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][2][4] [14]), .ZN(n_17_34_130));
   AOI22_X1 i_17_34_146 (.A1(\buffer[9][2][4] [14]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][2][4] [14]), .ZN(n_17_34_131));
   AOI22_X1 i_17_34_147 (.A1(\buffer[14][2][4] [14]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][2][4] [14]), .ZN(n_17_34_132));
   AOI22_X1 i_17_34_148 (.A1(\buffer[11][2][4] [14]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][2][4] [14]), .ZN(n_17_34_133));
   AOI22_X1 i_17_34_149 (.A1(\buffer[13][2][4] [14]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][2][4] [14]), .ZN(n_17_34_134));
   NAND2_X1 i_17_34_150 (.A1(n_17_34_137), .A2(n_17_34_135), .ZN(
      \output_filter[2][4] [15]));
   AOI221_X1 i_17_34_151 (.A(n_17_34_136), .B1(n_31), .B2(\buffer[3][2][4] [15]), 
      .C1(\buffer[14][2][4] [15]), .C2(n_19), .ZN(n_17_34_135));
   NAND3_X1 i_17_34_152 (.A1(n_17_34_143), .A2(n_17_34_141), .A3(n_17_34_139), 
      .ZN(n_17_34_136));
   AOI221_X1 i_17_34_153 (.A(n_17_34_138), .B1(n_16), .B2(\buffer[8][2][4] [15]), 
      .C1(\buffer[13][2][4] [15]), .C2(n_26), .ZN(n_17_34_137));
   NAND3_X1 i_17_34_154 (.A1(n_17_34_144), .A2(n_17_34_142), .A3(n_17_34_140), 
      .ZN(n_17_34_138));
   AOI22_X1 i_17_34_155 (.A1(\buffer[11][2][4] [15]), .A2(n_17), .B1(n_24), 
      .B2(\buffer[2][2][4] [15]), .ZN(n_17_34_139));
   AOI22_X1 i_17_34_156 (.A1(\buffer[10][2][4] [15]), .A2(n_21), .B1(n_23), 
      .B2(\buffer[1][2][4] [15]), .ZN(n_17_34_140));
   AOI22_X1 i_17_34_157 (.A1(\buffer[6][2][4] [15]), .A2(n_28), .B1(n_18), 
      .B2(\buffer[5][2][4] [15]), .ZN(n_17_34_141));
   AOI22_X1 i_17_34_158 (.A1(\buffer[9][2][4] [15]), .A2(n_20), .B1(n_30), 
      .B2(\buffer[4][2][4] [15]), .ZN(n_17_34_142));
   AOI22_X1 i_17_34_159 (.A1(\buffer[7][2][4] [15]), .A2(n_29), .B1(n_25), 
      .B2(\buffer[0][2][4] [15]), .ZN(n_17_34_143));
   AOI22_X1 i_17_34_160 (.A1(\buffer[15][2][4] [15]), .A2(n_22), .B1(n_27), 
      .B2(\buffer[12][2][4] [15]), .ZN(n_17_34_144));
   NAND4_X1 i_27_27_0 (.A1(n_27_27_8), .A2(n_27_27_6), .A3(n_27_27_4), .A4(
      n_27_27_0), .ZN(\output_filter[1][2] [0]));
   AOI221_X1 i_27_27_1 (.A(n_27_27_1), .B1(n_25), .B2(\buffer[0][1][2] [0]), 
      .C1(\buffer[12][1][2] [0]), .C2(n_27), .ZN(n_27_27_0));
   NAND4_X1 i_27_27_2 (.A1(n_27_27_7), .A2(n_27_27_5), .A3(n_27_27_3), .A4(
      n_27_27_2), .ZN(n_27_27_1));
   AOI22_X1 i_27_27_3 (.A1(\buffer[15][1][2] [0]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][2] [0]), .ZN(n_27_27_2));
   AOI22_X1 i_27_27_4 (.A1(\buffer[10][1][2] [0]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][2] [0]), .ZN(n_27_27_3));
   AOI22_X1 i_27_27_5 (.A1(\buffer[6][1][2] [0]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][1][2] [0]), .ZN(n_27_27_4));
   AOI22_X1 i_27_27_6 (.A1(\buffer[9][1][2] [0]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][1][2] [0]), .ZN(n_27_27_5));
   AOI22_X1 i_27_27_7 (.A1(\buffer[14][1][2] [0]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][2] [0]), .ZN(n_27_27_6));
   AOI22_X1 i_27_27_8 (.A1(\buffer[11][1][2] [0]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][2] [0]), .ZN(n_27_27_7));
   AOI22_X1 i_27_27_9 (.A1(\buffer[13][1][2] [0]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][2] [0]), .ZN(n_27_27_8));
   NAND4_X1 i_27_27_10 (.A1(n_27_27_17), .A2(n_27_27_15), .A3(n_27_27_13), 
      .A4(n_27_27_9), .ZN(\output_filter[1][2] [1]));
   AOI221_X1 i_27_27_11 (.A(n_27_27_10), .B1(n_25), .B2(\buffer[0][1][2] [1]), 
      .C1(\buffer[12][1][2] [1]), .C2(n_27), .ZN(n_27_27_9));
   NAND4_X1 i_27_27_12 (.A1(n_27_27_16), .A2(n_27_27_14), .A3(n_27_27_12), 
      .A4(n_27_27_11), .ZN(n_27_27_10));
   AOI22_X1 i_27_27_13 (.A1(\buffer[15][1][2] [1]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][2] [1]), .ZN(n_27_27_11));
   AOI22_X1 i_27_27_14 (.A1(\buffer[10][1][2] [1]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][2] [1]), .ZN(n_27_27_12));
   AOI22_X1 i_27_27_15 (.A1(\buffer[6][1][2] [1]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][2] [1]), .ZN(n_27_27_13));
   AOI22_X1 i_27_27_16 (.A1(\buffer[9][1][2] [1]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][2] [1]), .ZN(n_27_27_14));
   AOI22_X1 i_27_27_17 (.A1(\buffer[14][1][2] [1]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][2] [1]), .ZN(n_27_27_15));
   AOI22_X1 i_27_27_18 (.A1(\buffer[11][1][2] [1]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][2] [1]), .ZN(n_27_27_16));
   AOI22_X1 i_27_27_19 (.A1(\buffer[13][1][2] [1]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][2] [1]), .ZN(n_27_27_17));
   NAND4_X1 i_27_27_20 (.A1(n_27_27_26), .A2(n_27_27_24), .A3(n_27_27_22), 
      .A4(n_27_27_18), .ZN(\output_filter[1][2] [2]));
   AOI221_X1 i_27_27_21 (.A(n_27_27_19), .B1(n_25), .B2(\buffer[0][1][2] [2]), 
      .C1(\buffer[12][1][2] [2]), .C2(n_27), .ZN(n_27_27_18));
   NAND4_X1 i_27_27_22 (.A1(n_27_27_25), .A2(n_27_27_23), .A3(n_27_27_21), 
      .A4(n_27_27_20), .ZN(n_27_27_19));
   AOI22_X1 i_27_27_23 (.A1(\buffer[15][1][2] [2]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][2] [2]), .ZN(n_27_27_20));
   AOI22_X1 i_27_27_24 (.A1(\buffer[10][1][2] [2]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][2] [2]), .ZN(n_27_27_21));
   AOI22_X1 i_27_27_25 (.A1(\buffer[6][1][2] [2]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][2] [2]), .ZN(n_27_27_22));
   AOI22_X1 i_27_27_26 (.A1(\buffer[9][1][2] [2]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][2] [2]), .ZN(n_27_27_23));
   AOI22_X1 i_27_27_27 (.A1(\buffer[14][1][2] [2]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][2] [2]), .ZN(n_27_27_24));
   AOI22_X1 i_27_27_28 (.A1(\buffer[11][1][2] [2]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][2] [2]), .ZN(n_27_27_25));
   AOI22_X1 i_27_27_29 (.A1(\buffer[13][1][2] [2]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][2] [2]), .ZN(n_27_27_26));
   NAND4_X1 i_27_27_30 (.A1(n_27_27_35), .A2(n_27_27_33), .A3(n_27_27_31), 
      .A4(n_27_27_27), .ZN(\output_filter[1][2] [3]));
   AOI221_X1 i_27_27_31 (.A(n_27_27_28), .B1(n_25), .B2(\buffer[0][1][2] [3]), 
      .C1(\buffer[12][1][2] [3]), .C2(n_27), .ZN(n_27_27_27));
   NAND4_X1 i_27_27_32 (.A1(n_27_27_34), .A2(n_27_27_32), .A3(n_27_27_30), 
      .A4(n_27_27_29), .ZN(n_27_27_28));
   AOI22_X1 i_27_27_33 (.A1(\buffer[15][1][2] [3]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][2] [3]), .ZN(n_27_27_29));
   AOI22_X1 i_27_27_34 (.A1(\buffer[10][1][2] [3]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][2] [3]), .ZN(n_27_27_30));
   AOI22_X1 i_27_27_35 (.A1(\buffer[6][1][2] [3]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][2] [3]), .ZN(n_27_27_31));
   AOI22_X1 i_27_27_36 (.A1(\buffer[9][1][2] [3]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][2] [3]), .ZN(n_27_27_32));
   AOI22_X1 i_27_27_37 (.A1(\buffer[14][1][2] [3]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][2] [3]), .ZN(n_27_27_33));
   AOI22_X1 i_27_27_38 (.A1(\buffer[11][1][2] [3]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][2] [3]), .ZN(n_27_27_34));
   AOI22_X1 i_27_27_39 (.A1(\buffer[13][1][2] [3]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][2] [3]), .ZN(n_27_27_35));
   NAND4_X1 i_27_27_40 (.A1(n_27_27_44), .A2(n_27_27_42), .A3(n_27_27_40), 
      .A4(n_27_27_36), .ZN(\output_filter[1][2] [4]));
   AOI221_X1 i_27_27_41 (.A(n_27_27_37), .B1(n_25), .B2(\buffer[0][1][2] [4]), 
      .C1(\buffer[12][1][2] [4]), .C2(n_27), .ZN(n_27_27_36));
   NAND4_X1 i_27_27_42 (.A1(n_27_27_43), .A2(n_27_27_41), .A3(n_27_27_39), 
      .A4(n_27_27_38), .ZN(n_27_27_37));
   AOI22_X1 i_27_27_43 (.A1(\buffer[15][1][2] [4]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][2] [4]), .ZN(n_27_27_38));
   AOI22_X1 i_27_27_44 (.A1(\buffer[10][1][2] [4]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][2] [4]), .ZN(n_27_27_39));
   AOI22_X1 i_27_27_45 (.A1(\buffer[6][1][2] [4]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][2] [4]), .ZN(n_27_27_40));
   AOI22_X1 i_27_27_46 (.A1(\buffer[9][1][2] [4]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][1][2] [4]), .ZN(n_27_27_41));
   AOI22_X1 i_27_27_47 (.A1(\buffer[14][1][2] [4]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][2] [4]), .ZN(n_27_27_42));
   AOI22_X1 i_27_27_48 (.A1(\buffer[11][1][2] [4]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][2] [4]), .ZN(n_27_27_43));
   AOI22_X1 i_27_27_49 (.A1(\buffer[13][1][2] [4]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][1][2] [4]), .ZN(n_27_27_44));
   NAND4_X1 i_27_27_50 (.A1(n_27_27_53), .A2(n_27_27_51), .A3(n_27_27_49), 
      .A4(n_27_27_45), .ZN(\output_filter[1][2] [5]));
   AOI221_X1 i_27_27_51 (.A(n_27_27_46), .B1(n_25), .B2(\buffer[0][1][2] [5]), 
      .C1(\buffer[12][1][2] [5]), .C2(n_27), .ZN(n_27_27_45));
   NAND4_X1 i_27_27_52 (.A1(n_27_27_52), .A2(n_27_27_50), .A3(n_27_27_48), 
      .A4(n_27_27_47), .ZN(n_27_27_46));
   AOI22_X1 i_27_27_53 (.A1(\buffer[15][1][2] [5]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][2] [5]), .ZN(n_27_27_47));
   AOI22_X1 i_27_27_54 (.A1(\buffer[10][1][2] [5]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][2] [5]), .ZN(n_27_27_48));
   AOI22_X1 i_27_27_55 (.A1(\buffer[6][1][2] [5]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][2] [5]), .ZN(n_27_27_49));
   AOI22_X1 i_27_27_56 (.A1(\buffer[9][1][2] [5]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][2] [5]), .ZN(n_27_27_50));
   AOI22_X1 i_27_27_57 (.A1(\buffer[14][1][2] [5]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][2] [5]), .ZN(n_27_27_51));
   AOI22_X1 i_27_27_58 (.A1(\buffer[11][1][2] [5]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][2] [5]), .ZN(n_27_27_52));
   AOI22_X1 i_27_27_59 (.A1(\buffer[13][1][2] [5]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][2] [5]), .ZN(n_27_27_53));
   NAND4_X1 i_27_27_60 (.A1(n_27_27_62), .A2(n_27_27_60), .A3(n_27_27_58), 
      .A4(n_27_27_54), .ZN(\output_filter[1][2] [6]));
   AOI221_X1 i_27_27_61 (.A(n_27_27_55), .B1(n_25), .B2(\buffer[0][1][2] [6]), 
      .C1(\buffer[12][1][2] [6]), .C2(n_27), .ZN(n_27_27_54));
   NAND4_X1 i_27_27_62 (.A1(n_27_27_61), .A2(n_27_27_59), .A3(n_27_27_57), 
      .A4(n_27_27_56), .ZN(n_27_27_55));
   AOI22_X1 i_27_27_63 (.A1(\buffer[15][1][2] [6]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][2] [6]), .ZN(n_27_27_56));
   AOI22_X1 i_27_27_64 (.A1(\buffer[10][1][2] [6]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][2] [6]), .ZN(n_27_27_57));
   AOI22_X1 i_27_27_65 (.A1(\buffer[6][1][2] [6]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][2] [6]), .ZN(n_27_27_58));
   AOI22_X1 i_27_27_66 (.A1(\buffer[9][1][2] [6]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][2] [6]), .ZN(n_27_27_59));
   AOI22_X1 i_27_27_67 (.A1(\buffer[14][1][2] [6]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][2] [6]), .ZN(n_27_27_60));
   AOI22_X1 i_27_27_68 (.A1(\buffer[11][1][2] [6]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][2] [6]), .ZN(n_27_27_61));
   AOI22_X1 i_27_27_69 (.A1(\buffer[13][1][2] [6]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][2] [6]), .ZN(n_27_27_62));
   NAND4_X1 i_27_27_70 (.A1(n_27_27_71), .A2(n_27_27_69), .A3(n_27_27_67), 
      .A4(n_27_27_63), .ZN(\output_filter[1][2] [7]));
   AOI221_X1 i_27_27_71 (.A(n_27_27_64), .B1(n_25), .B2(\buffer[0][1][2] [7]), 
      .C1(\buffer[12][1][2] [7]), .C2(n_27), .ZN(n_27_27_63));
   NAND4_X1 i_27_27_72 (.A1(n_27_27_70), .A2(n_27_27_68), .A3(n_27_27_66), 
      .A4(n_27_27_65), .ZN(n_27_27_64));
   AOI22_X1 i_27_27_73 (.A1(\buffer[15][1][2] [7]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][2] [7]), .ZN(n_27_27_65));
   AOI22_X1 i_27_27_74 (.A1(\buffer[10][1][2] [7]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][2] [7]), .ZN(n_27_27_66));
   AOI22_X1 i_27_27_75 (.A1(\buffer[6][1][2] [7]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][2] [7]), .ZN(n_27_27_67));
   AOI22_X1 i_27_27_76 (.A1(\buffer[9][1][2] [7]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][1][2] [7]), .ZN(n_27_27_68));
   AOI22_X1 i_27_27_77 (.A1(\buffer[14][1][2] [7]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][2] [7]), .ZN(n_27_27_69));
   AOI22_X1 i_27_27_78 (.A1(\buffer[11][1][2] [7]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][2] [7]), .ZN(n_27_27_70));
   AOI22_X1 i_27_27_79 (.A1(\buffer[13][1][2] [7]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][1][2] [7]), .ZN(n_27_27_71));
   NAND4_X1 i_27_27_80 (.A1(n_27_27_80), .A2(n_27_27_78), .A3(n_27_27_76), 
      .A4(n_27_27_72), .ZN(\output_filter[1][2] [8]));
   AOI221_X1 i_27_27_81 (.A(n_27_27_73), .B1(n_25), .B2(\buffer[0][1][2] [8]), 
      .C1(\buffer[12][1][2] [8]), .C2(n_27), .ZN(n_27_27_72));
   NAND4_X1 i_27_27_82 (.A1(n_27_27_79), .A2(n_27_27_77), .A3(n_27_27_75), 
      .A4(n_27_27_74), .ZN(n_27_27_73));
   AOI22_X1 i_27_27_83 (.A1(\buffer[15][1][2] [8]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][2] [8]), .ZN(n_27_27_74));
   AOI22_X1 i_27_27_84 (.A1(\buffer[10][1][2] [8]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][2] [8]), .ZN(n_27_27_75));
   AOI22_X1 i_27_27_85 (.A1(\buffer[6][1][2] [8]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][2] [8]), .ZN(n_27_27_76));
   AOI22_X1 i_27_27_86 (.A1(\buffer[9][1][2] [8]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][2] [8]), .ZN(n_27_27_77));
   AOI22_X1 i_27_27_87 (.A1(\buffer[14][1][2] [8]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][2] [8]), .ZN(n_27_27_78));
   AOI22_X1 i_27_27_88 (.A1(\buffer[11][1][2] [8]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][2] [8]), .ZN(n_27_27_79));
   AOI22_X1 i_27_27_89 (.A1(\buffer[13][1][2] [8]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][2] [8]), .ZN(n_27_27_80));
   NAND4_X1 i_27_27_90 (.A1(n_27_27_89), .A2(n_27_27_87), .A3(n_27_27_85), 
      .A4(n_27_27_81), .ZN(\output_filter[1][2] [9]));
   AOI221_X1 i_27_27_91 (.A(n_27_27_82), .B1(n_25), .B2(\buffer[0][1][2] [9]), 
      .C1(\buffer[12][1][2] [9]), .C2(n_27), .ZN(n_27_27_81));
   NAND4_X1 i_27_27_92 (.A1(n_27_27_88), .A2(n_27_27_86), .A3(n_27_27_84), 
      .A4(n_27_27_83), .ZN(n_27_27_82));
   AOI22_X1 i_27_27_93 (.A1(\buffer[15][1][2] [9]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][2] [9]), .ZN(n_27_27_83));
   AOI22_X1 i_27_27_94 (.A1(\buffer[10][1][2] [9]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][2] [9]), .ZN(n_27_27_84));
   AOI22_X1 i_27_27_95 (.A1(\buffer[6][1][2] [9]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][2] [9]), .ZN(n_27_27_85));
   AOI22_X1 i_27_27_96 (.A1(\buffer[9][1][2] [9]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][1][2] [9]), .ZN(n_27_27_86));
   AOI22_X1 i_27_27_97 (.A1(\buffer[14][1][2] [9]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][2] [9]), .ZN(n_27_27_87));
   AOI22_X1 i_27_27_98 (.A1(\buffer[11][1][2] [9]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][2] [9]), .ZN(n_27_27_88));
   AOI22_X1 i_27_27_99 (.A1(\buffer[13][1][2] [9]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][1][2] [9]), .ZN(n_27_27_89));
   NAND4_X1 i_27_27_100 (.A1(n_27_27_98), .A2(n_27_27_96), .A3(n_27_27_94), 
      .A4(n_27_27_90), .ZN(\output_filter[1][2] [10]));
   AOI221_X1 i_27_27_101 (.A(n_27_27_91), .B1(n_25), .B2(\buffer[0][1][2] [10]), 
      .C1(\buffer[12][1][2] [10]), .C2(n_27), .ZN(n_27_27_90));
   NAND4_X1 i_27_27_102 (.A1(n_27_27_97), .A2(n_27_27_95), .A3(n_27_27_93), 
      .A4(n_27_27_92), .ZN(n_27_27_91));
   AOI22_X1 i_27_27_103 (.A1(\buffer[15][1][2] [10]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][2] [10]), .ZN(n_27_27_92));
   AOI22_X1 i_27_27_104 (.A1(\buffer[10][1][2] [10]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][2] [10]), .ZN(n_27_27_93));
   AOI22_X1 i_27_27_105 (.A1(\buffer[6][1][2] [10]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][2] [10]), .ZN(n_27_27_94));
   AOI22_X1 i_27_27_106 (.A1(\buffer[9][1][2] [10]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][2] [10]), .ZN(n_27_27_95));
   AOI22_X1 i_27_27_107 (.A1(\buffer[14][1][2] [10]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][2] [10]), .ZN(n_27_27_96));
   AOI22_X1 i_27_27_108 (.A1(\buffer[11][1][2] [10]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][2] [10]), .ZN(n_27_27_97));
   AOI22_X1 i_27_27_109 (.A1(\buffer[13][1][2] [10]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][2] [10]), .ZN(n_27_27_98));
   NAND4_X1 i_27_27_110 (.A1(n_27_27_107), .A2(n_27_27_105), .A3(n_27_27_103), 
      .A4(n_27_27_99), .ZN(\output_filter[1][2] [11]));
   AOI221_X1 i_27_27_111 (.A(n_27_27_100), .B1(n_25), .B2(\buffer[0][1][2] [11]), 
      .C1(\buffer[12][1][2] [11]), .C2(n_27), .ZN(n_27_27_99));
   NAND4_X1 i_27_27_112 (.A1(n_27_27_106), .A2(n_27_27_104), .A3(n_27_27_102), 
      .A4(n_27_27_101), .ZN(n_27_27_100));
   AOI22_X1 i_27_27_113 (.A1(\buffer[15][1][2] [11]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][2] [11]), .ZN(n_27_27_101));
   AOI22_X1 i_27_27_114 (.A1(\buffer[10][1][2] [11]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][2] [11]), .ZN(n_27_27_102));
   AOI22_X1 i_27_27_115 (.A1(\buffer[6][1][2] [11]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][2] [11]), .ZN(n_27_27_103));
   AOI22_X1 i_27_27_116 (.A1(\buffer[9][1][2] [11]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][1][2] [11]), .ZN(n_27_27_104));
   AOI22_X1 i_27_27_117 (.A1(\buffer[14][1][2] [11]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][2] [11]), .ZN(n_27_27_105));
   AOI22_X1 i_27_27_118 (.A1(\buffer[11][1][2] [11]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][2] [11]), .ZN(n_27_27_106));
   AOI22_X1 i_27_27_119 (.A1(\buffer[13][1][2] [11]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][1][2] [11]), .ZN(n_27_27_107));
   NAND4_X1 i_27_27_120 (.A1(n_27_27_116), .A2(n_27_27_114), .A3(n_27_27_112), 
      .A4(n_27_27_108), .ZN(\output_filter[1][2] [12]));
   AOI221_X1 i_27_27_121 (.A(n_27_27_109), .B1(n_25), .B2(\buffer[0][1][2] [12]), 
      .C1(\buffer[12][1][2] [12]), .C2(n_27), .ZN(n_27_27_108));
   NAND4_X1 i_27_27_122 (.A1(n_27_27_115), .A2(n_27_27_113), .A3(n_27_27_111), 
      .A4(n_27_27_110), .ZN(n_27_27_109));
   AOI22_X1 i_27_27_123 (.A1(\buffer[15][1][2] [12]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][2] [12]), .ZN(n_27_27_110));
   AOI22_X1 i_27_27_124 (.A1(\buffer[10][1][2] [12]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][2] [12]), .ZN(n_27_27_111));
   AOI22_X1 i_27_27_125 (.A1(\buffer[6][1][2] [12]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][2] [12]), .ZN(n_27_27_112));
   AOI22_X1 i_27_27_126 (.A1(\buffer[9][1][2] [12]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][2] [12]), .ZN(n_27_27_113));
   AOI22_X1 i_27_27_127 (.A1(\buffer[14][1][2] [12]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][2] [12]), .ZN(n_27_27_114));
   AOI22_X1 i_27_27_128 (.A1(\buffer[11][1][2] [12]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][2] [12]), .ZN(n_27_27_115));
   AOI22_X1 i_27_27_129 (.A1(\buffer[13][1][2] [12]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][2] [12]), .ZN(n_27_27_116));
   NAND4_X1 i_27_27_130 (.A1(n_27_27_125), .A2(n_27_27_123), .A3(n_27_27_121), 
      .A4(n_27_27_117), .ZN(\output_filter[1][2] [13]));
   AOI221_X1 i_27_27_131 (.A(n_27_27_118), .B1(n_25), .B2(\buffer[0][1][2] [13]), 
      .C1(\buffer[12][1][2] [13]), .C2(n_27), .ZN(n_27_27_117));
   NAND4_X1 i_27_27_132 (.A1(n_27_27_124), .A2(n_27_27_122), .A3(n_27_27_120), 
      .A4(n_27_27_119), .ZN(n_27_27_118));
   AOI22_X1 i_27_27_133 (.A1(\buffer[15][1][2] [13]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][2] [13]), .ZN(n_27_27_119));
   AOI22_X1 i_27_27_134 (.A1(\buffer[10][1][2] [13]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][2] [13]), .ZN(n_27_27_120));
   AOI22_X1 i_27_27_135 (.A1(\buffer[6][1][2] [13]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][2] [13]), .ZN(n_27_27_121));
   AOI22_X1 i_27_27_136 (.A1(\buffer[9][1][2] [13]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][1][2] [13]), .ZN(n_27_27_122));
   AOI22_X1 i_27_27_137 (.A1(\buffer[14][1][2] [13]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][2] [13]), .ZN(n_27_27_123));
   AOI22_X1 i_27_27_138 (.A1(\buffer[11][1][2] [13]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][2] [13]), .ZN(n_27_27_124));
   AOI22_X1 i_27_27_139 (.A1(\buffer[13][1][2] [13]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][1][2] [13]), .ZN(n_27_27_125));
   NAND4_X1 i_27_27_140 (.A1(n_27_27_134), .A2(n_27_27_132), .A3(n_27_27_130), 
      .A4(n_27_27_126), .ZN(\output_filter[1][2] [14]));
   AOI221_X1 i_27_27_141 (.A(n_27_27_127), .B1(n_25), .B2(\buffer[0][1][2] [14]), 
      .C1(\buffer[12][1][2] [14]), .C2(n_27), .ZN(n_27_27_126));
   NAND4_X1 i_27_27_142 (.A1(n_27_27_133), .A2(n_27_27_131), .A3(n_27_27_129), 
      .A4(n_27_27_128), .ZN(n_27_27_127));
   AOI22_X1 i_27_27_143 (.A1(\buffer[15][1][2] [14]), .A2(n_22), .B1(n_16), 
      .B2(\buffer[8][1][2] [14]), .ZN(n_27_27_128));
   AOI22_X1 i_27_27_144 (.A1(\buffer[10][1][2] [14]), .A2(n_21), .B1(n_29), 
      .B2(\buffer[7][1][2] [14]), .ZN(n_27_27_129));
   AOI22_X1 i_27_27_145 (.A1(\buffer[6][1][2] [14]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][2] [14]), .ZN(n_27_27_130));
   AOI22_X1 i_27_27_146 (.A1(\buffer[9][1][2] [14]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][2] [14]), .ZN(n_27_27_131));
   AOI22_X1 i_27_27_147 (.A1(\buffer[14][1][2] [14]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][2] [14]), .ZN(n_27_27_132));
   AOI22_X1 i_27_27_148 (.A1(\buffer[11][1][2] [14]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][2] [14]), .ZN(n_27_27_133));
   AOI22_X1 i_27_27_149 (.A1(\buffer[13][1][2] [14]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][2] [14]), .ZN(n_27_27_134));
   NAND2_X1 i_27_27_150 (.A1(n_27_27_137), .A2(n_27_27_135), .ZN(
      \output_filter[1][2] [15]));
   AOI221_X1 i_27_27_151 (.A(n_27_27_136), .B1(n_31), .B2(\buffer[3][1][2] [15]), 
      .C1(\buffer[14][1][2] [15]), .C2(n_19), .ZN(n_27_27_135));
   NAND3_X1 i_27_27_152 (.A1(n_27_27_143), .A2(n_27_27_141), .A3(n_27_27_139), 
      .ZN(n_27_27_136));
   AOI221_X1 i_27_27_153 (.A(n_27_27_138), .B1(n_16), .B2(\buffer[8][1][2] [15]), 
      .C1(\buffer[13][1][2] [15]), .C2(n_26), .ZN(n_27_27_137));
   NAND3_X1 i_27_27_154 (.A1(n_27_27_144), .A2(n_27_27_142), .A3(n_27_27_140), 
      .ZN(n_27_27_138));
   AOI22_X1 i_27_27_155 (.A1(\buffer[11][1][2] [15]), .A2(n_17), .B1(n_24), 
      .B2(\buffer[2][1][2] [15]), .ZN(n_27_27_139));
   AOI22_X1 i_27_27_156 (.A1(\buffer[10][1][2] [15]), .A2(n_21), .B1(n_23), 
      .B2(\buffer[1][1][2] [15]), .ZN(n_27_27_140));
   AOI22_X1 i_27_27_157 (.A1(\buffer[6][1][2] [15]), .A2(n_28), .B1(n_18), 
      .B2(\buffer[5][1][2] [15]), .ZN(n_27_27_141));
   AOI22_X1 i_27_27_158 (.A1(\buffer[9][1][2] [15]), .A2(n_20), .B1(n_30), 
      .B2(\buffer[4][1][2] [15]), .ZN(n_27_27_142));
   AOI22_X1 i_27_27_159 (.A1(\buffer[7][1][2] [15]), .A2(n_29), .B1(n_25), 
      .B2(\buffer[0][1][2] [15]), .ZN(n_27_27_143));
   AOI22_X1 i_27_27_160 (.A1(\buffer[15][1][2] [15]), .A2(n_22), .B1(n_27), 
      .B2(\buffer[12][1][2] [15]), .ZN(n_27_27_144));
   NAND4_X1 i_26_26_0 (.A1(n_26_26_8), .A2(n_26_26_6), .A3(n_26_26_4), .A4(
      n_26_26_0), .ZN(\output_filter[1][1] [0]));
   AOI221_X1 i_26_26_1 (.A(n_26_26_1), .B1(n_25), .B2(\buffer[0][1][1] [0]), 
      .C1(\buffer[12][1][1] [0]), .C2(n_27), .ZN(n_26_26_0));
   NAND4_X1 i_26_26_2 (.A1(n_26_26_7), .A2(n_26_26_5), .A3(n_26_26_3), .A4(
      n_26_26_2), .ZN(n_26_26_1));
   AOI22_X1 i_26_26_3 (.A1(\buffer[15][1][1] [0]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][1] [0]), .ZN(n_26_26_2));
   AOI22_X1 i_26_26_4 (.A1(\buffer[10][1][1] [0]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][1] [0]), .ZN(n_26_26_3));
   AOI22_X1 i_26_26_5 (.A1(\buffer[6][1][1] [0]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][1][1] [0]), .ZN(n_26_26_4));
   AOI22_X1 i_26_26_6 (.A1(\buffer[9][1][1] [0]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][1][1] [0]), .ZN(n_26_26_5));
   AOI22_X1 i_26_26_7 (.A1(\buffer[14][1][1] [0]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][1] [0]), .ZN(n_26_26_6));
   AOI22_X1 i_26_26_8 (.A1(\buffer[11][1][1] [0]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][1] [0]), .ZN(n_26_26_7));
   AOI22_X1 i_26_26_9 (.A1(\buffer[13][1][1] [0]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][1] [0]), .ZN(n_26_26_8));
   NAND4_X1 i_26_26_10 (.A1(n_26_26_17), .A2(n_26_26_15), .A3(n_26_26_13), 
      .A4(n_26_26_9), .ZN(\output_filter[1][1] [1]));
   AOI221_X1 i_26_26_11 (.A(n_26_26_10), .B1(n_25), .B2(\buffer[0][1][1] [1]), 
      .C1(\buffer[12][1][1] [1]), .C2(n_27), .ZN(n_26_26_9));
   NAND4_X1 i_26_26_12 (.A1(n_26_26_16), .A2(n_26_26_14), .A3(n_26_26_12), 
      .A4(n_26_26_11), .ZN(n_26_26_10));
   AOI22_X1 i_26_26_13 (.A1(\buffer[15][1][1] [1]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][1] [1]), .ZN(n_26_26_11));
   AOI22_X1 i_26_26_14 (.A1(\buffer[10][1][1] [1]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][1] [1]), .ZN(n_26_26_12));
   AOI22_X1 i_26_26_15 (.A1(\buffer[6][1][1] [1]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][1] [1]), .ZN(n_26_26_13));
   AOI22_X1 i_26_26_16 (.A1(\buffer[9][1][1] [1]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][1] [1]), .ZN(n_26_26_14));
   AOI22_X1 i_26_26_17 (.A1(\buffer[14][1][1] [1]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][1] [1]), .ZN(n_26_26_15));
   AOI22_X1 i_26_26_18 (.A1(\buffer[11][1][1] [1]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][1] [1]), .ZN(n_26_26_16));
   AOI22_X1 i_26_26_19 (.A1(\buffer[13][1][1] [1]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][1] [1]), .ZN(n_26_26_17));
   NAND4_X1 i_26_26_20 (.A1(n_26_26_26), .A2(n_26_26_24), .A3(n_26_26_22), 
      .A4(n_26_26_18), .ZN(\output_filter[1][1] [2]));
   AOI221_X1 i_26_26_21 (.A(n_26_26_19), .B1(n_25), .B2(\buffer[0][1][1] [2]), 
      .C1(\buffer[12][1][1] [2]), .C2(n_27), .ZN(n_26_26_18));
   NAND4_X1 i_26_26_22 (.A1(n_26_26_25), .A2(n_26_26_23), .A3(n_26_26_21), 
      .A4(n_26_26_20), .ZN(n_26_26_19));
   AOI22_X1 i_26_26_23 (.A1(\buffer[15][1][1] [2]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][1] [2]), .ZN(n_26_26_20));
   AOI22_X1 i_26_26_24 (.A1(\buffer[10][1][1] [2]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][1] [2]), .ZN(n_26_26_21));
   AOI22_X1 i_26_26_25 (.A1(\buffer[6][1][1] [2]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][1] [2]), .ZN(n_26_26_22));
   AOI22_X1 i_26_26_26 (.A1(\buffer[9][1][1] [2]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][1] [2]), .ZN(n_26_26_23));
   AOI22_X1 i_26_26_27 (.A1(\buffer[14][1][1] [2]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][1] [2]), .ZN(n_26_26_24));
   AOI22_X1 i_26_26_28 (.A1(\buffer[11][1][1] [2]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][1] [2]), .ZN(n_26_26_25));
   AOI22_X1 i_26_26_29 (.A1(\buffer[13][1][1] [2]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][1] [2]), .ZN(n_26_26_26));
   NAND4_X1 i_26_26_30 (.A1(n_26_26_35), .A2(n_26_26_33), .A3(n_26_26_31), 
      .A4(n_26_26_27), .ZN(\output_filter[1][1] [3]));
   AOI221_X1 i_26_26_31 (.A(n_26_26_28), .B1(n_25), .B2(\buffer[0][1][1] [3]), 
      .C1(\buffer[12][1][1] [3]), .C2(n_27), .ZN(n_26_26_27));
   NAND4_X1 i_26_26_32 (.A1(n_26_26_34), .A2(n_26_26_32), .A3(n_26_26_30), 
      .A4(n_26_26_29), .ZN(n_26_26_28));
   AOI22_X1 i_26_26_33 (.A1(\buffer[15][1][1] [3]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][1] [3]), .ZN(n_26_26_29));
   AOI22_X1 i_26_26_34 (.A1(\buffer[10][1][1] [3]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][1] [3]), .ZN(n_26_26_30));
   AOI22_X1 i_26_26_35 (.A1(\buffer[6][1][1] [3]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][1] [3]), .ZN(n_26_26_31));
   AOI22_X1 i_26_26_36 (.A1(\buffer[9][1][1] [3]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][1] [3]), .ZN(n_26_26_32));
   AOI22_X1 i_26_26_37 (.A1(\buffer[14][1][1] [3]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][1] [3]), .ZN(n_26_26_33));
   AOI22_X1 i_26_26_38 (.A1(\buffer[11][1][1] [3]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][1] [3]), .ZN(n_26_26_34));
   AOI22_X1 i_26_26_39 (.A1(\buffer[13][1][1] [3]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][1] [3]), .ZN(n_26_26_35));
   NAND4_X1 i_26_26_40 (.A1(n_26_26_44), .A2(n_26_26_42), .A3(n_26_26_40), 
      .A4(n_26_26_36), .ZN(\output_filter[1][1] [4]));
   AOI221_X1 i_26_26_41 (.A(n_26_26_37), .B1(n_25), .B2(\buffer[0][1][1] [4]), 
      .C1(\buffer[12][1][1] [4]), .C2(n_27), .ZN(n_26_26_36));
   NAND4_X1 i_26_26_42 (.A1(n_26_26_43), .A2(n_26_26_41), .A3(n_26_26_39), 
      .A4(n_26_26_38), .ZN(n_26_26_37));
   AOI22_X1 i_26_26_43 (.A1(\buffer[15][1][1] [4]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][1] [4]), .ZN(n_26_26_38));
   AOI22_X1 i_26_26_44 (.A1(\buffer[10][1][1] [4]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][1] [4]), .ZN(n_26_26_39));
   AOI22_X1 i_26_26_45 (.A1(\buffer[6][1][1] [4]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][1] [4]), .ZN(n_26_26_40));
   AOI22_X1 i_26_26_46 (.A1(\buffer[9][1][1] [4]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][1][1] [4]), .ZN(n_26_26_41));
   AOI22_X1 i_26_26_47 (.A1(\buffer[14][1][1] [4]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][1] [4]), .ZN(n_26_26_42));
   AOI22_X1 i_26_26_48 (.A1(\buffer[11][1][1] [4]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][1] [4]), .ZN(n_26_26_43));
   AOI22_X1 i_26_26_49 (.A1(\buffer[13][1][1] [4]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][1][1] [4]), .ZN(n_26_26_44));
   NAND4_X1 i_26_26_50 (.A1(n_26_26_53), .A2(n_26_26_51), .A3(n_26_26_49), 
      .A4(n_26_26_45), .ZN(\output_filter[1][1] [5]));
   AOI221_X1 i_26_26_51 (.A(n_26_26_46), .B1(n_25), .B2(\buffer[0][1][1] [5]), 
      .C1(\buffer[12][1][1] [5]), .C2(n_27), .ZN(n_26_26_45));
   NAND4_X1 i_26_26_52 (.A1(n_26_26_52), .A2(n_26_26_50), .A3(n_26_26_48), 
      .A4(n_26_26_47), .ZN(n_26_26_46));
   AOI22_X1 i_26_26_53 (.A1(\buffer[15][1][1] [5]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][1] [5]), .ZN(n_26_26_47));
   AOI22_X1 i_26_26_54 (.A1(\buffer[10][1][1] [5]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][1] [5]), .ZN(n_26_26_48));
   AOI22_X1 i_26_26_55 (.A1(\buffer[6][1][1] [5]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][1] [5]), .ZN(n_26_26_49));
   AOI22_X1 i_26_26_56 (.A1(\buffer[9][1][1] [5]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][1] [5]), .ZN(n_26_26_50));
   AOI22_X1 i_26_26_57 (.A1(\buffer[14][1][1] [5]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][1] [5]), .ZN(n_26_26_51));
   AOI22_X1 i_26_26_58 (.A1(\buffer[11][1][1] [5]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][1] [5]), .ZN(n_26_26_52));
   AOI22_X1 i_26_26_59 (.A1(\buffer[13][1][1] [5]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][1] [5]), .ZN(n_26_26_53));
   NAND4_X1 i_26_26_60 (.A1(n_26_26_62), .A2(n_26_26_60), .A3(n_26_26_58), 
      .A4(n_26_26_54), .ZN(\output_filter[1][1] [6]));
   AOI221_X1 i_26_26_61 (.A(n_26_26_55), .B1(n_25), .B2(\buffer[0][1][1] [6]), 
      .C1(\buffer[12][1][1] [6]), .C2(n_27), .ZN(n_26_26_54));
   NAND4_X1 i_26_26_62 (.A1(n_26_26_61), .A2(n_26_26_59), .A3(n_26_26_57), 
      .A4(n_26_26_56), .ZN(n_26_26_55));
   AOI22_X1 i_26_26_63 (.A1(\buffer[15][1][1] [6]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][1] [6]), .ZN(n_26_26_56));
   AOI22_X1 i_26_26_64 (.A1(\buffer[10][1][1] [6]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][1] [6]), .ZN(n_26_26_57));
   AOI22_X1 i_26_26_65 (.A1(\buffer[6][1][1] [6]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][1] [6]), .ZN(n_26_26_58));
   AOI22_X1 i_26_26_66 (.A1(\buffer[9][1][1] [6]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][1] [6]), .ZN(n_26_26_59));
   AOI22_X1 i_26_26_67 (.A1(\buffer[14][1][1] [6]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][1] [6]), .ZN(n_26_26_60));
   AOI22_X1 i_26_26_68 (.A1(\buffer[11][1][1] [6]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][1] [6]), .ZN(n_26_26_61));
   AOI22_X1 i_26_26_69 (.A1(\buffer[13][1][1] [6]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][1] [6]), .ZN(n_26_26_62));
   NAND4_X1 i_26_26_70 (.A1(n_26_26_71), .A2(n_26_26_69), .A3(n_26_26_67), 
      .A4(n_26_26_63), .ZN(\output_filter[1][1] [7]));
   AOI221_X1 i_26_26_71 (.A(n_26_26_64), .B1(n_25), .B2(\buffer[0][1][1] [7]), 
      .C1(\buffer[12][1][1] [7]), .C2(n_27), .ZN(n_26_26_63));
   NAND4_X1 i_26_26_72 (.A1(n_26_26_70), .A2(n_26_26_68), .A3(n_26_26_66), 
      .A4(n_26_26_65), .ZN(n_26_26_64));
   AOI22_X1 i_26_26_73 (.A1(\buffer[15][1][1] [7]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][1] [7]), .ZN(n_26_26_65));
   AOI22_X1 i_26_26_74 (.A1(\buffer[10][1][1] [7]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][1] [7]), .ZN(n_26_26_66));
   AOI22_X1 i_26_26_75 (.A1(\buffer[6][1][1] [7]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][1] [7]), .ZN(n_26_26_67));
   AOI22_X1 i_26_26_76 (.A1(\buffer[9][1][1] [7]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][1][1] [7]), .ZN(n_26_26_68));
   AOI22_X1 i_26_26_77 (.A1(\buffer[14][1][1] [7]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][1] [7]), .ZN(n_26_26_69));
   AOI22_X1 i_26_26_78 (.A1(\buffer[11][1][1] [7]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][1] [7]), .ZN(n_26_26_70));
   AOI22_X1 i_26_26_79 (.A1(\buffer[13][1][1] [7]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][1][1] [7]), .ZN(n_26_26_71));
   NAND4_X1 i_26_26_80 (.A1(n_26_26_80), .A2(n_26_26_78), .A3(n_26_26_76), 
      .A4(n_26_26_72), .ZN(\output_filter[1][1] [8]));
   AOI221_X1 i_26_26_81 (.A(n_26_26_73), .B1(n_25), .B2(\buffer[0][1][1] [8]), 
      .C1(\buffer[12][1][1] [8]), .C2(n_27), .ZN(n_26_26_72));
   NAND4_X1 i_26_26_82 (.A1(n_26_26_79), .A2(n_26_26_77), .A3(n_26_26_75), 
      .A4(n_26_26_74), .ZN(n_26_26_73));
   AOI22_X1 i_26_26_83 (.A1(\buffer[15][1][1] [8]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][1] [8]), .ZN(n_26_26_74));
   AOI22_X1 i_26_26_84 (.A1(\buffer[10][1][1] [8]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][1] [8]), .ZN(n_26_26_75));
   AOI22_X1 i_26_26_85 (.A1(\buffer[6][1][1] [8]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][1] [8]), .ZN(n_26_26_76));
   AOI22_X1 i_26_26_86 (.A1(\buffer[9][1][1] [8]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][1] [8]), .ZN(n_26_26_77));
   AOI22_X1 i_26_26_87 (.A1(\buffer[14][1][1] [8]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][1] [8]), .ZN(n_26_26_78));
   AOI22_X1 i_26_26_88 (.A1(\buffer[11][1][1] [8]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][1] [8]), .ZN(n_26_26_79));
   AOI22_X1 i_26_26_89 (.A1(\buffer[13][1][1] [8]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][1] [8]), .ZN(n_26_26_80));
   NAND4_X1 i_26_26_90 (.A1(n_26_26_89), .A2(n_26_26_87), .A3(n_26_26_85), 
      .A4(n_26_26_81), .ZN(\output_filter[1][1] [9]));
   AOI221_X1 i_26_26_91 (.A(n_26_26_82), .B1(n_25), .B2(\buffer[0][1][1] [9]), 
      .C1(\buffer[12][1][1] [9]), .C2(n_27), .ZN(n_26_26_81));
   NAND4_X1 i_26_26_92 (.A1(n_26_26_88), .A2(n_26_26_86), .A3(n_26_26_84), 
      .A4(n_26_26_83), .ZN(n_26_26_82));
   AOI22_X1 i_26_26_93 (.A1(\buffer[15][1][1] [9]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][1] [9]), .ZN(n_26_26_83));
   AOI22_X1 i_26_26_94 (.A1(\buffer[10][1][1] [9]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][1] [9]), .ZN(n_26_26_84));
   AOI22_X1 i_26_26_95 (.A1(\buffer[6][1][1] [9]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][1] [9]), .ZN(n_26_26_85));
   AOI22_X1 i_26_26_96 (.A1(\buffer[9][1][1] [9]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][1][1] [9]), .ZN(n_26_26_86));
   AOI22_X1 i_26_26_97 (.A1(\buffer[14][1][1] [9]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][1] [9]), .ZN(n_26_26_87));
   AOI22_X1 i_26_26_98 (.A1(\buffer[11][1][1] [9]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][1] [9]), .ZN(n_26_26_88));
   AOI22_X1 i_26_26_99 (.A1(\buffer[13][1][1] [9]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][1][1] [9]), .ZN(n_26_26_89));
   NAND4_X1 i_26_26_100 (.A1(n_26_26_98), .A2(n_26_26_96), .A3(n_26_26_94), 
      .A4(n_26_26_90), .ZN(\output_filter[1][1] [10]));
   AOI221_X1 i_26_26_101 (.A(n_26_26_91), .B1(n_25), .B2(\buffer[0][1][1] [10]), 
      .C1(\buffer[12][1][1] [10]), .C2(n_27), .ZN(n_26_26_90));
   NAND4_X1 i_26_26_102 (.A1(n_26_26_97), .A2(n_26_26_95), .A3(n_26_26_93), 
      .A4(n_26_26_92), .ZN(n_26_26_91));
   AOI22_X1 i_26_26_103 (.A1(\buffer[15][1][1] [10]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][1] [10]), .ZN(n_26_26_92));
   AOI22_X1 i_26_26_104 (.A1(\buffer[10][1][1] [10]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][1] [10]), .ZN(n_26_26_93));
   AOI22_X1 i_26_26_105 (.A1(\buffer[6][1][1] [10]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][1] [10]), .ZN(n_26_26_94));
   AOI22_X1 i_26_26_106 (.A1(\buffer[9][1][1] [10]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][1] [10]), .ZN(n_26_26_95));
   AOI22_X1 i_26_26_107 (.A1(\buffer[14][1][1] [10]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][1] [10]), .ZN(n_26_26_96));
   AOI22_X1 i_26_26_108 (.A1(\buffer[11][1][1] [10]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][1] [10]), .ZN(n_26_26_97));
   AOI22_X1 i_26_26_109 (.A1(\buffer[13][1][1] [10]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][1] [10]), .ZN(n_26_26_98));
   NAND4_X1 i_26_26_110 (.A1(n_26_26_107), .A2(n_26_26_105), .A3(n_26_26_103), 
      .A4(n_26_26_99), .ZN(\output_filter[1][1] [11]));
   AOI221_X1 i_26_26_111 (.A(n_26_26_100), .B1(n_25), .B2(\buffer[0][1][1] [11]), 
      .C1(\buffer[12][1][1] [11]), .C2(n_27), .ZN(n_26_26_99));
   NAND4_X1 i_26_26_112 (.A1(n_26_26_106), .A2(n_26_26_104), .A3(n_26_26_102), 
      .A4(n_26_26_101), .ZN(n_26_26_100));
   AOI22_X1 i_26_26_113 (.A1(\buffer[15][1][1] [11]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][1] [11]), .ZN(n_26_26_101));
   AOI22_X1 i_26_26_114 (.A1(\buffer[10][1][1] [11]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][1] [11]), .ZN(n_26_26_102));
   AOI22_X1 i_26_26_115 (.A1(\buffer[6][1][1] [11]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][1] [11]), .ZN(n_26_26_103));
   AOI22_X1 i_26_26_116 (.A1(\buffer[9][1][1] [11]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][1][1] [11]), .ZN(n_26_26_104));
   AOI22_X1 i_26_26_117 (.A1(\buffer[14][1][1] [11]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][1] [11]), .ZN(n_26_26_105));
   AOI22_X1 i_26_26_118 (.A1(\buffer[11][1][1] [11]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][1] [11]), .ZN(n_26_26_106));
   AOI22_X1 i_26_26_119 (.A1(\buffer[13][1][1] [11]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][1][1] [11]), .ZN(n_26_26_107));
   NAND4_X1 i_26_26_120 (.A1(n_26_26_116), .A2(n_26_26_114), .A3(n_26_26_112), 
      .A4(n_26_26_108), .ZN(\output_filter[1][1] [12]));
   AOI221_X1 i_26_26_121 (.A(n_26_26_109), .B1(n_25), .B2(\buffer[0][1][1] [12]), 
      .C1(\buffer[12][1][1] [12]), .C2(n_27), .ZN(n_26_26_108));
   NAND4_X1 i_26_26_122 (.A1(n_26_26_115), .A2(n_26_26_113), .A3(n_26_26_111), 
      .A4(n_26_26_110), .ZN(n_26_26_109));
   AOI22_X1 i_26_26_123 (.A1(\buffer[15][1][1] [12]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][1] [12]), .ZN(n_26_26_110));
   AOI22_X1 i_26_26_124 (.A1(\buffer[10][1][1] [12]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][1] [12]), .ZN(n_26_26_111));
   AOI22_X1 i_26_26_125 (.A1(\buffer[6][1][1] [12]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][1] [12]), .ZN(n_26_26_112));
   AOI22_X1 i_26_26_126 (.A1(\buffer[9][1][1] [12]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][1] [12]), .ZN(n_26_26_113));
   AOI22_X1 i_26_26_127 (.A1(\buffer[14][1][1] [12]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][1] [12]), .ZN(n_26_26_114));
   AOI22_X1 i_26_26_128 (.A1(\buffer[11][1][1] [12]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][1] [12]), .ZN(n_26_26_115));
   AOI22_X1 i_26_26_129 (.A1(\buffer[13][1][1] [12]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][1] [12]), .ZN(n_26_26_116));
   NAND4_X1 i_26_26_130 (.A1(n_26_26_125), .A2(n_26_26_123), .A3(n_26_26_121), 
      .A4(n_26_26_117), .ZN(\output_filter[1][1] [13]));
   AOI221_X1 i_26_26_131 (.A(n_26_26_118), .B1(n_25), .B2(\buffer[0][1][1] [13]), 
      .C1(\buffer[12][1][1] [13]), .C2(n_27), .ZN(n_26_26_117));
   NAND4_X1 i_26_26_132 (.A1(n_26_26_124), .A2(n_26_26_122), .A3(n_26_26_120), 
      .A4(n_26_26_119), .ZN(n_26_26_118));
   AOI22_X1 i_26_26_133 (.A1(\buffer[15][1][1] [13]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][1] [13]), .ZN(n_26_26_119));
   AOI22_X1 i_26_26_134 (.A1(\buffer[10][1][1] [13]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][1] [13]), .ZN(n_26_26_120));
   AOI22_X1 i_26_26_135 (.A1(\buffer[6][1][1] [13]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][1] [13]), .ZN(n_26_26_121));
   AOI22_X1 i_26_26_136 (.A1(\buffer[9][1][1] [13]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][1][1] [13]), .ZN(n_26_26_122));
   AOI22_X1 i_26_26_137 (.A1(\buffer[14][1][1] [13]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][1] [13]), .ZN(n_26_26_123));
   AOI22_X1 i_26_26_138 (.A1(\buffer[11][1][1] [13]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][1] [13]), .ZN(n_26_26_124));
   AOI22_X1 i_26_26_139 (.A1(\buffer[13][1][1] [13]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][1][1] [13]), .ZN(n_26_26_125));
   NAND4_X1 i_26_26_140 (.A1(n_26_26_134), .A2(n_26_26_132), .A3(n_26_26_130), 
      .A4(n_26_26_126), .ZN(\output_filter[1][1] [14]));
   AOI221_X1 i_26_26_141 (.A(n_26_26_127), .B1(n_25), .B2(\buffer[0][1][1] [14]), 
      .C1(\buffer[12][1][1] [14]), .C2(n_27), .ZN(n_26_26_126));
   NAND4_X1 i_26_26_142 (.A1(n_26_26_133), .A2(n_26_26_131), .A3(n_26_26_129), 
      .A4(n_26_26_128), .ZN(n_26_26_127));
   AOI22_X1 i_26_26_143 (.A1(\buffer[15][1][1] [14]), .A2(n_22), .B1(n_16), 
      .B2(\buffer[8][1][1] [14]), .ZN(n_26_26_128));
   AOI22_X1 i_26_26_144 (.A1(\buffer[10][1][1] [14]), .A2(n_21), .B1(n_29), 
      .B2(\buffer[7][1][1] [14]), .ZN(n_26_26_129));
   AOI22_X1 i_26_26_145 (.A1(\buffer[6][1][1] [14]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][1] [14]), .ZN(n_26_26_130));
   AOI22_X1 i_26_26_146 (.A1(\buffer[9][1][1] [14]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][1] [14]), .ZN(n_26_26_131));
   AOI22_X1 i_26_26_147 (.A1(\buffer[14][1][1] [14]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][1] [14]), .ZN(n_26_26_132));
   AOI22_X1 i_26_26_148 (.A1(\buffer[11][1][1] [14]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][1] [14]), .ZN(n_26_26_133));
   AOI22_X1 i_26_26_149 (.A1(\buffer[13][1][1] [14]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][1] [14]), .ZN(n_26_26_134));
   NAND2_X1 i_26_26_150 (.A1(n_26_26_137), .A2(n_26_26_135), .ZN(
      \output_filter[1][1] [15]));
   AOI221_X1 i_26_26_151 (.A(n_26_26_136), .B1(n_31), .B2(\buffer[3][1][1] [15]), 
      .C1(\buffer[14][1][1] [15]), .C2(n_19), .ZN(n_26_26_135));
   NAND3_X1 i_26_26_152 (.A1(n_26_26_143), .A2(n_26_26_141), .A3(n_26_26_139), 
      .ZN(n_26_26_136));
   AOI221_X1 i_26_26_153 (.A(n_26_26_138), .B1(n_16), .B2(\buffer[8][1][1] [15]), 
      .C1(\buffer[13][1][1] [15]), .C2(n_26), .ZN(n_26_26_137));
   NAND3_X1 i_26_26_154 (.A1(n_26_26_144), .A2(n_26_26_142), .A3(n_26_26_140), 
      .ZN(n_26_26_138));
   AOI22_X1 i_26_26_155 (.A1(\buffer[11][1][1] [15]), .A2(n_17), .B1(n_24), 
      .B2(\buffer[2][1][1] [15]), .ZN(n_26_26_139));
   AOI22_X1 i_26_26_156 (.A1(\buffer[10][1][1] [15]), .A2(n_21), .B1(n_23), 
      .B2(\buffer[1][1][1] [15]), .ZN(n_26_26_140));
   AOI22_X1 i_26_26_157 (.A1(\buffer[6][1][1] [15]), .A2(n_28), .B1(n_18), 
      .B2(\buffer[5][1][1] [15]), .ZN(n_26_26_141));
   AOI22_X1 i_26_26_158 (.A1(\buffer[9][1][1] [15]), .A2(n_20), .B1(n_30), 
      .B2(\buffer[4][1][1] [15]), .ZN(n_26_26_142));
   AOI22_X1 i_26_26_159 (.A1(\buffer[7][1][1] [15]), .A2(n_29), .B1(n_25), 
      .B2(\buffer[0][1][1] [15]), .ZN(n_26_26_143));
   AOI22_X1 i_26_26_160 (.A1(\buffer[15][1][1] [15]), .A2(n_22), .B1(n_27), 
      .B2(\buffer[12][1][1] [15]), .ZN(n_26_26_144));
   NAND4_X1 i_25_25_0 (.A1(n_25_25_8), .A2(n_25_25_6), .A3(n_25_25_4), .A4(
      n_25_25_0), .ZN(\output_filter[1][0] [0]));
   AOI221_X1 i_25_25_1 (.A(n_25_25_1), .B1(n_25), .B2(\buffer[0][1][0] [0]), 
      .C1(\buffer[12][1][0] [0]), .C2(n_27), .ZN(n_25_25_0));
   NAND4_X1 i_25_25_2 (.A1(n_25_25_7), .A2(n_25_25_5), .A3(n_25_25_3), .A4(
      n_25_25_2), .ZN(n_25_25_1));
   AOI22_X1 i_25_25_3 (.A1(\buffer[15][1][0] [0]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][0] [0]), .ZN(n_25_25_2));
   AOI22_X1 i_25_25_4 (.A1(\buffer[10][1][0] [0]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][0] [0]), .ZN(n_25_25_3));
   AOI22_X1 i_25_25_5 (.A1(\buffer[6][1][0] [0]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][1][0] [0]), .ZN(n_25_25_4));
   AOI22_X1 i_25_25_6 (.A1(\buffer[9][1][0] [0]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][1][0] [0]), .ZN(n_25_25_5));
   AOI22_X1 i_25_25_7 (.A1(\buffer[14][1][0] [0]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][0] [0]), .ZN(n_25_25_6));
   AOI22_X1 i_25_25_8 (.A1(\buffer[11][1][0] [0]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][0] [0]), .ZN(n_25_25_7));
   AOI22_X1 i_25_25_9 (.A1(\buffer[13][1][0] [0]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][0] [0]), .ZN(n_25_25_8));
   NAND4_X1 i_25_25_10 (.A1(n_25_25_17), .A2(n_25_25_15), .A3(n_25_25_13), 
      .A4(n_25_25_9), .ZN(\output_filter[1][0] [1]));
   AOI221_X1 i_25_25_11 (.A(n_25_25_10), .B1(n_25), .B2(\buffer[0][1][0] [1]), 
      .C1(\buffer[12][1][0] [1]), .C2(n_27), .ZN(n_25_25_9));
   NAND4_X1 i_25_25_12 (.A1(n_25_25_16), .A2(n_25_25_14), .A3(n_25_25_12), 
      .A4(n_25_25_11), .ZN(n_25_25_10));
   AOI22_X1 i_25_25_13 (.A1(\buffer[15][1][0] [1]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][0] [1]), .ZN(n_25_25_11));
   AOI22_X1 i_25_25_14 (.A1(\buffer[10][1][0] [1]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][0] [1]), .ZN(n_25_25_12));
   AOI22_X1 i_25_25_15 (.A1(\buffer[6][1][0] [1]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][0] [1]), .ZN(n_25_25_13));
   AOI22_X1 i_25_25_16 (.A1(\buffer[9][1][0] [1]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][0] [1]), .ZN(n_25_25_14));
   AOI22_X1 i_25_25_17 (.A1(\buffer[14][1][0] [1]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][0] [1]), .ZN(n_25_25_15));
   AOI22_X1 i_25_25_18 (.A1(\buffer[11][1][0] [1]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][0] [1]), .ZN(n_25_25_16));
   AOI22_X1 i_25_25_19 (.A1(\buffer[13][1][0] [1]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][0] [1]), .ZN(n_25_25_17));
   NAND4_X1 i_25_25_20 (.A1(n_25_25_26), .A2(n_25_25_24), .A3(n_25_25_22), 
      .A4(n_25_25_18), .ZN(\output_filter[1][0] [2]));
   AOI221_X1 i_25_25_21 (.A(n_25_25_19), .B1(n_25), .B2(\buffer[0][1][0] [2]), 
      .C1(\buffer[12][1][0] [2]), .C2(n_27), .ZN(n_25_25_18));
   NAND4_X1 i_25_25_22 (.A1(n_25_25_25), .A2(n_25_25_23), .A3(n_25_25_21), 
      .A4(n_25_25_20), .ZN(n_25_25_19));
   AOI22_X1 i_25_25_23 (.A1(\buffer[15][1][0] [2]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][0] [2]), .ZN(n_25_25_20));
   AOI22_X1 i_25_25_24 (.A1(\buffer[10][1][0] [2]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][0] [2]), .ZN(n_25_25_21));
   AOI22_X1 i_25_25_25 (.A1(\buffer[6][1][0] [2]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][0] [2]), .ZN(n_25_25_22));
   AOI22_X1 i_25_25_26 (.A1(\buffer[9][1][0] [2]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][0] [2]), .ZN(n_25_25_23));
   AOI22_X1 i_25_25_27 (.A1(\buffer[14][1][0] [2]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][0] [2]), .ZN(n_25_25_24));
   AOI22_X1 i_25_25_28 (.A1(\buffer[11][1][0] [2]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][0] [2]), .ZN(n_25_25_25));
   AOI22_X1 i_25_25_29 (.A1(\buffer[13][1][0] [2]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][0] [2]), .ZN(n_25_25_26));
   NAND4_X1 i_25_25_30 (.A1(n_25_25_35), .A2(n_25_25_33), .A3(n_25_25_31), 
      .A4(n_25_25_27), .ZN(\output_filter[1][0] [3]));
   AOI221_X1 i_25_25_31 (.A(n_25_25_28), .B1(n_25), .B2(\buffer[0][1][0] [3]), 
      .C1(\buffer[12][1][0] [3]), .C2(n_27), .ZN(n_25_25_27));
   NAND4_X1 i_25_25_32 (.A1(n_25_25_34), .A2(n_25_25_32), .A3(n_25_25_30), 
      .A4(n_25_25_29), .ZN(n_25_25_28));
   AOI22_X1 i_25_25_33 (.A1(\buffer[15][1][0] [3]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][0] [3]), .ZN(n_25_25_29));
   AOI22_X1 i_25_25_34 (.A1(\buffer[10][1][0] [3]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][0] [3]), .ZN(n_25_25_30));
   AOI22_X1 i_25_25_35 (.A1(\buffer[6][1][0] [3]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][0] [3]), .ZN(n_25_25_31));
   AOI22_X1 i_25_25_36 (.A1(\buffer[9][1][0] [3]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][0] [3]), .ZN(n_25_25_32));
   AOI22_X1 i_25_25_37 (.A1(\buffer[14][1][0] [3]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][0] [3]), .ZN(n_25_25_33));
   AOI22_X1 i_25_25_38 (.A1(\buffer[11][1][0] [3]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][0] [3]), .ZN(n_25_25_34));
   AOI22_X1 i_25_25_39 (.A1(\buffer[13][1][0] [3]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][0] [3]), .ZN(n_25_25_35));
   NAND4_X1 i_25_25_40 (.A1(n_25_25_44), .A2(n_25_25_42), .A3(n_25_25_40), 
      .A4(n_25_25_36), .ZN(\output_filter[1][0] [4]));
   AOI221_X1 i_25_25_41 (.A(n_25_25_37), .B1(n_25), .B2(\buffer[0][1][0] [4]), 
      .C1(\buffer[12][1][0] [4]), .C2(n_27), .ZN(n_25_25_36));
   NAND4_X1 i_25_25_42 (.A1(n_25_25_43), .A2(n_25_25_41), .A3(n_25_25_39), 
      .A4(n_25_25_38), .ZN(n_25_25_37));
   AOI22_X1 i_25_25_43 (.A1(\buffer[15][1][0] [4]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][0] [4]), .ZN(n_25_25_38));
   AOI22_X1 i_25_25_44 (.A1(\buffer[10][1][0] [4]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][0] [4]), .ZN(n_25_25_39));
   AOI22_X1 i_25_25_45 (.A1(\buffer[6][1][0] [4]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][0] [4]), .ZN(n_25_25_40));
   AOI22_X1 i_25_25_46 (.A1(\buffer[9][1][0] [4]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][1][0] [4]), .ZN(n_25_25_41));
   AOI22_X1 i_25_25_47 (.A1(\buffer[14][1][0] [4]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][0] [4]), .ZN(n_25_25_42));
   AOI22_X1 i_25_25_48 (.A1(\buffer[11][1][0] [4]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][0] [4]), .ZN(n_25_25_43));
   AOI22_X1 i_25_25_49 (.A1(\buffer[13][1][0] [4]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][1][0] [4]), .ZN(n_25_25_44));
   NAND4_X1 i_25_25_50 (.A1(n_25_25_53), .A2(n_25_25_51), .A3(n_25_25_49), 
      .A4(n_25_25_45), .ZN(\output_filter[1][0] [5]));
   AOI221_X1 i_25_25_51 (.A(n_25_25_46), .B1(n_25), .B2(\buffer[0][1][0] [5]), 
      .C1(\buffer[12][1][0] [5]), .C2(n_27), .ZN(n_25_25_45));
   NAND4_X1 i_25_25_52 (.A1(n_25_25_52), .A2(n_25_25_50), .A3(n_25_25_48), 
      .A4(n_25_25_47), .ZN(n_25_25_46));
   AOI22_X1 i_25_25_53 (.A1(\buffer[15][1][0] [5]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][0] [5]), .ZN(n_25_25_47));
   AOI22_X1 i_25_25_54 (.A1(\buffer[10][1][0] [5]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][0] [5]), .ZN(n_25_25_48));
   AOI22_X1 i_25_25_55 (.A1(\buffer[6][1][0] [5]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][0] [5]), .ZN(n_25_25_49));
   AOI22_X1 i_25_25_56 (.A1(\buffer[9][1][0] [5]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][0] [5]), .ZN(n_25_25_50));
   AOI22_X1 i_25_25_57 (.A1(\buffer[14][1][0] [5]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][0] [5]), .ZN(n_25_25_51));
   AOI22_X1 i_25_25_58 (.A1(\buffer[11][1][0] [5]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][0] [5]), .ZN(n_25_25_52));
   AOI22_X1 i_25_25_59 (.A1(\buffer[13][1][0] [5]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][0] [5]), .ZN(n_25_25_53));
   NAND4_X1 i_25_25_60 (.A1(n_25_25_62), .A2(n_25_25_60), .A3(n_25_25_58), 
      .A4(n_25_25_54), .ZN(\output_filter[1][0] [6]));
   AOI221_X1 i_25_25_61 (.A(n_25_25_55), .B1(n_25), .B2(\buffer[0][1][0] [6]), 
      .C1(\buffer[12][1][0] [6]), .C2(n_27), .ZN(n_25_25_54));
   NAND4_X1 i_25_25_62 (.A1(n_25_25_61), .A2(n_25_25_59), .A3(n_25_25_57), 
      .A4(n_25_25_56), .ZN(n_25_25_55));
   AOI22_X1 i_25_25_63 (.A1(\buffer[15][1][0] [6]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][0] [6]), .ZN(n_25_25_56));
   AOI22_X1 i_25_25_64 (.A1(\buffer[10][1][0] [6]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][0] [6]), .ZN(n_25_25_57));
   AOI22_X1 i_25_25_65 (.A1(\buffer[6][1][0] [6]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][0] [6]), .ZN(n_25_25_58));
   AOI22_X1 i_25_25_66 (.A1(\buffer[9][1][0] [6]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][0] [6]), .ZN(n_25_25_59));
   AOI22_X1 i_25_25_67 (.A1(\buffer[14][1][0] [6]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][0] [6]), .ZN(n_25_25_60));
   AOI22_X1 i_25_25_68 (.A1(\buffer[11][1][0] [6]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][0] [6]), .ZN(n_25_25_61));
   AOI22_X1 i_25_25_69 (.A1(\buffer[13][1][0] [6]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][0] [6]), .ZN(n_25_25_62));
   NAND4_X1 i_25_25_70 (.A1(n_25_25_71), .A2(n_25_25_69), .A3(n_25_25_67), 
      .A4(n_25_25_63), .ZN(\output_filter[1][0] [7]));
   AOI221_X1 i_25_25_71 (.A(n_25_25_64), .B1(n_25), .B2(\buffer[0][1][0] [7]), 
      .C1(\buffer[12][1][0] [7]), .C2(n_27), .ZN(n_25_25_63));
   NAND4_X1 i_25_25_72 (.A1(n_25_25_70), .A2(n_25_25_68), .A3(n_25_25_66), 
      .A4(n_25_25_65), .ZN(n_25_25_64));
   AOI22_X1 i_25_25_73 (.A1(\buffer[15][1][0] [7]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][0] [7]), .ZN(n_25_25_65));
   AOI22_X1 i_25_25_74 (.A1(\buffer[10][1][0] [7]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][0] [7]), .ZN(n_25_25_66));
   AOI22_X1 i_25_25_75 (.A1(\buffer[6][1][0] [7]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][0] [7]), .ZN(n_25_25_67));
   AOI22_X1 i_25_25_76 (.A1(\buffer[9][1][0] [7]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][1][0] [7]), .ZN(n_25_25_68));
   AOI22_X1 i_25_25_77 (.A1(\buffer[14][1][0] [7]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][0] [7]), .ZN(n_25_25_69));
   AOI22_X1 i_25_25_78 (.A1(\buffer[11][1][0] [7]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][0] [7]), .ZN(n_25_25_70));
   AOI22_X1 i_25_25_79 (.A1(\buffer[13][1][0] [7]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][1][0] [7]), .ZN(n_25_25_71));
   NAND4_X1 i_25_25_80 (.A1(n_25_25_80), .A2(n_25_25_78), .A3(n_25_25_76), 
      .A4(n_25_25_72), .ZN(\output_filter[1][0] [8]));
   AOI221_X1 i_25_25_81 (.A(n_25_25_73), .B1(n_25), .B2(\buffer[0][1][0] [8]), 
      .C1(\buffer[12][1][0] [8]), .C2(n_27), .ZN(n_25_25_72));
   NAND4_X1 i_25_25_82 (.A1(n_25_25_79), .A2(n_25_25_77), .A3(n_25_25_75), 
      .A4(n_25_25_74), .ZN(n_25_25_73));
   AOI22_X1 i_25_25_83 (.A1(\buffer[15][1][0] [8]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][0] [8]), .ZN(n_25_25_74));
   AOI22_X1 i_25_25_84 (.A1(\buffer[10][1][0] [8]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][0] [8]), .ZN(n_25_25_75));
   AOI22_X1 i_25_25_85 (.A1(\buffer[6][1][0] [8]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][0] [8]), .ZN(n_25_25_76));
   AOI22_X1 i_25_25_86 (.A1(\buffer[9][1][0] [8]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][0] [8]), .ZN(n_25_25_77));
   AOI22_X1 i_25_25_87 (.A1(\buffer[14][1][0] [8]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][0] [8]), .ZN(n_25_25_78));
   AOI22_X1 i_25_25_88 (.A1(\buffer[11][1][0] [8]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][0] [8]), .ZN(n_25_25_79));
   AOI22_X1 i_25_25_89 (.A1(\buffer[13][1][0] [8]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][0] [8]), .ZN(n_25_25_80));
   NAND4_X1 i_25_25_90 (.A1(n_25_25_89), .A2(n_25_25_87), .A3(n_25_25_85), 
      .A4(n_25_25_81), .ZN(\output_filter[1][0] [9]));
   AOI221_X1 i_25_25_91 (.A(n_25_25_82), .B1(n_25), .B2(\buffer[0][1][0] [9]), 
      .C1(\buffer[12][1][0] [9]), .C2(n_27), .ZN(n_25_25_81));
   NAND4_X1 i_25_25_92 (.A1(n_25_25_88), .A2(n_25_25_86), .A3(n_25_25_84), 
      .A4(n_25_25_83), .ZN(n_25_25_82));
   AOI22_X1 i_25_25_93 (.A1(\buffer[15][1][0] [9]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][0] [9]), .ZN(n_25_25_83));
   AOI22_X1 i_25_25_94 (.A1(\buffer[10][1][0] [9]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][0] [9]), .ZN(n_25_25_84));
   AOI22_X1 i_25_25_95 (.A1(\buffer[6][1][0] [9]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][0] [9]), .ZN(n_25_25_85));
   AOI22_X1 i_25_25_96 (.A1(\buffer[9][1][0] [9]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][1][0] [9]), .ZN(n_25_25_86));
   AOI22_X1 i_25_25_97 (.A1(\buffer[14][1][0] [9]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][0] [9]), .ZN(n_25_25_87));
   AOI22_X1 i_25_25_98 (.A1(\buffer[11][1][0] [9]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][0] [9]), .ZN(n_25_25_88));
   AOI22_X1 i_25_25_99 (.A1(\buffer[13][1][0] [9]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][1][0] [9]), .ZN(n_25_25_89));
   NAND4_X1 i_25_25_100 (.A1(n_25_25_98), .A2(n_25_25_96), .A3(n_25_25_94), 
      .A4(n_25_25_90), .ZN(\output_filter[1][0] [10]));
   AOI221_X1 i_25_25_101 (.A(n_25_25_91), .B1(n_25), .B2(\buffer[0][1][0] [10]), 
      .C1(\buffer[12][1][0] [10]), .C2(n_27), .ZN(n_25_25_90));
   NAND4_X1 i_25_25_102 (.A1(n_25_25_97), .A2(n_25_25_95), .A3(n_25_25_93), 
      .A4(n_25_25_92), .ZN(n_25_25_91));
   AOI22_X1 i_25_25_103 (.A1(\buffer[15][1][0] [10]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][0] [10]), .ZN(n_25_25_92));
   AOI22_X1 i_25_25_104 (.A1(\buffer[10][1][0] [10]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][0] [10]), .ZN(n_25_25_93));
   AOI22_X1 i_25_25_105 (.A1(\buffer[6][1][0] [10]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][0] [10]), .ZN(n_25_25_94));
   AOI22_X1 i_25_25_106 (.A1(\buffer[9][1][0] [10]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][0] [10]), .ZN(n_25_25_95));
   AOI22_X1 i_25_25_107 (.A1(\buffer[14][1][0] [10]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][0] [10]), .ZN(n_25_25_96));
   AOI22_X1 i_25_25_108 (.A1(\buffer[11][1][0] [10]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][0] [10]), .ZN(n_25_25_97));
   AOI22_X1 i_25_25_109 (.A1(\buffer[13][1][0] [10]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][0] [10]), .ZN(n_25_25_98));
   NAND4_X1 i_25_25_110 (.A1(n_25_25_107), .A2(n_25_25_105), .A3(n_25_25_103), 
      .A4(n_25_25_99), .ZN(\output_filter[1][0] [11]));
   AOI221_X1 i_25_25_111 (.A(n_25_25_100), .B1(n_25), .B2(\buffer[0][1][0] [11]), 
      .C1(\buffer[12][1][0] [11]), .C2(n_27), .ZN(n_25_25_99));
   NAND4_X1 i_25_25_112 (.A1(n_25_25_106), .A2(n_25_25_104), .A3(n_25_25_102), 
      .A4(n_25_25_101), .ZN(n_25_25_100));
   AOI22_X1 i_25_25_113 (.A1(\buffer[15][1][0] [11]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][0] [11]), .ZN(n_25_25_101));
   AOI22_X1 i_25_25_114 (.A1(\buffer[10][1][0] [11]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][0] [11]), .ZN(n_25_25_102));
   AOI22_X1 i_25_25_115 (.A1(\buffer[6][1][0] [11]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][0] [11]), .ZN(n_25_25_103));
   AOI22_X1 i_25_25_116 (.A1(\buffer[9][1][0] [11]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][1][0] [11]), .ZN(n_25_25_104));
   AOI22_X1 i_25_25_117 (.A1(\buffer[14][1][0] [11]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][0] [11]), .ZN(n_25_25_105));
   AOI22_X1 i_25_25_118 (.A1(\buffer[11][1][0] [11]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][0] [11]), .ZN(n_25_25_106));
   AOI22_X1 i_25_25_119 (.A1(\buffer[13][1][0] [11]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][1][0] [11]), .ZN(n_25_25_107));
   NAND4_X1 i_25_25_120 (.A1(n_25_25_116), .A2(n_25_25_114), .A3(n_25_25_112), 
      .A4(n_25_25_108), .ZN(\output_filter[1][0] [12]));
   AOI221_X1 i_25_25_121 (.A(n_25_25_109), .B1(n_25), .B2(\buffer[0][1][0] [12]), 
      .C1(\buffer[12][1][0] [12]), .C2(n_27), .ZN(n_25_25_108));
   NAND4_X1 i_25_25_122 (.A1(n_25_25_115), .A2(n_25_25_113), .A3(n_25_25_111), 
      .A4(n_25_25_110), .ZN(n_25_25_109));
   AOI22_X1 i_25_25_123 (.A1(\buffer[15][1][0] [12]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][0] [12]), .ZN(n_25_25_110));
   AOI22_X1 i_25_25_124 (.A1(\buffer[10][1][0] [12]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][0] [12]), .ZN(n_25_25_111));
   AOI22_X1 i_25_25_125 (.A1(\buffer[6][1][0] [12]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][0] [12]), .ZN(n_25_25_112));
   AOI22_X1 i_25_25_126 (.A1(\buffer[9][1][0] [12]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][0] [12]), .ZN(n_25_25_113));
   AOI22_X1 i_25_25_127 (.A1(\buffer[14][1][0] [12]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][0] [12]), .ZN(n_25_25_114));
   AOI22_X1 i_25_25_128 (.A1(\buffer[11][1][0] [12]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][0] [12]), .ZN(n_25_25_115));
   AOI22_X1 i_25_25_129 (.A1(\buffer[13][1][0] [12]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][0] [12]), .ZN(n_25_25_116));
   NAND4_X1 i_25_25_130 (.A1(n_25_25_125), .A2(n_25_25_123), .A3(n_25_25_121), 
      .A4(n_25_25_117), .ZN(\output_filter[1][0] [13]));
   AOI221_X1 i_25_25_131 (.A(n_25_25_118), .B1(n_25), .B2(\buffer[0][1][0] [13]), 
      .C1(\buffer[12][1][0] [13]), .C2(n_27), .ZN(n_25_25_117));
   NAND4_X1 i_25_25_132 (.A1(n_25_25_124), .A2(n_25_25_122), .A3(n_25_25_120), 
      .A4(n_25_25_119), .ZN(n_25_25_118));
   AOI22_X1 i_25_25_133 (.A1(\buffer[15][1][0] [13]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][1][0] [13]), .ZN(n_25_25_119));
   AOI22_X1 i_25_25_134 (.A1(\buffer[10][1][0] [13]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][1][0] [13]), .ZN(n_25_25_120));
   AOI22_X1 i_25_25_135 (.A1(\buffer[6][1][0] [13]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][0] [13]), .ZN(n_25_25_121));
   AOI22_X1 i_25_25_136 (.A1(\buffer[9][1][0] [13]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][1][0] [13]), .ZN(n_25_25_122));
   AOI22_X1 i_25_25_137 (.A1(\buffer[14][1][0] [13]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][0] [13]), .ZN(n_25_25_123));
   AOI22_X1 i_25_25_138 (.A1(\buffer[11][1][0] [13]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][0] [13]), .ZN(n_25_25_124));
   AOI22_X1 i_25_25_139 (.A1(\buffer[13][1][0] [13]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][1][0] [13]), .ZN(n_25_25_125));
   NAND4_X1 i_25_25_140 (.A1(n_25_25_134), .A2(n_25_25_132), .A3(n_25_25_130), 
      .A4(n_25_25_126), .ZN(\output_filter[1][0] [14]));
   AOI221_X1 i_25_25_141 (.A(n_25_25_127), .B1(n_25), .B2(\buffer[0][1][0] [14]), 
      .C1(\buffer[12][1][0] [14]), .C2(n_27), .ZN(n_25_25_126));
   NAND4_X1 i_25_25_142 (.A1(n_25_25_133), .A2(n_25_25_131), .A3(n_25_25_129), 
      .A4(n_25_25_128), .ZN(n_25_25_127));
   AOI22_X1 i_25_25_143 (.A1(\buffer[15][1][0] [14]), .A2(n_22), .B1(n_16), 
      .B2(\buffer[8][1][0] [14]), .ZN(n_25_25_128));
   AOI22_X1 i_25_25_144 (.A1(\buffer[10][1][0] [14]), .A2(n_21), .B1(n_29), 
      .B2(\buffer[7][1][0] [14]), .ZN(n_25_25_129));
   AOI22_X1 i_25_25_145 (.A1(\buffer[6][1][0] [14]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][1][0] [14]), .ZN(n_25_25_130));
   AOI22_X1 i_25_25_146 (.A1(\buffer[9][1][0] [14]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][1][0] [14]), .ZN(n_25_25_131));
   AOI22_X1 i_25_25_147 (.A1(\buffer[14][1][0] [14]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][1][0] [14]), .ZN(n_25_25_132));
   AOI22_X1 i_25_25_148 (.A1(\buffer[11][1][0] [14]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][1][0] [14]), .ZN(n_25_25_133));
   AOI22_X1 i_25_25_149 (.A1(\buffer[13][1][0] [14]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][1][0] [14]), .ZN(n_25_25_134));
   NAND2_X1 i_25_25_150 (.A1(n_25_25_137), .A2(n_25_25_135), .ZN(
      \output_filter[1][0] [15]));
   AOI221_X1 i_25_25_151 (.A(n_25_25_136), .B1(n_31), .B2(\buffer[3][1][0] [15]), 
      .C1(\buffer[14][1][0] [15]), .C2(n_19), .ZN(n_25_25_135));
   NAND3_X1 i_25_25_152 (.A1(n_25_25_143), .A2(n_25_25_141), .A3(n_25_25_139), 
      .ZN(n_25_25_136));
   AOI221_X1 i_25_25_153 (.A(n_25_25_138), .B1(n_16), .B2(\buffer[8][1][0] [15]), 
      .C1(\buffer[13][1][0] [15]), .C2(n_26), .ZN(n_25_25_137));
   NAND3_X1 i_25_25_154 (.A1(n_25_25_144), .A2(n_25_25_142), .A3(n_25_25_140), 
      .ZN(n_25_25_138));
   AOI22_X1 i_25_25_155 (.A1(\buffer[11][1][0] [15]), .A2(n_17), .B1(n_24), 
      .B2(\buffer[2][1][0] [15]), .ZN(n_25_25_139));
   AOI22_X1 i_25_25_156 (.A1(\buffer[10][1][0] [15]), .A2(n_21), .B1(n_23), 
      .B2(\buffer[1][1][0] [15]), .ZN(n_25_25_140));
   AOI22_X1 i_25_25_157 (.A1(\buffer[6][1][0] [15]), .A2(n_28), .B1(n_18), 
      .B2(\buffer[5][1][0] [15]), .ZN(n_25_25_141));
   AOI22_X1 i_25_25_158 (.A1(\buffer[9][1][0] [15]), .A2(n_20), .B1(n_30), 
      .B2(\buffer[4][1][0] [15]), .ZN(n_25_25_142));
   AOI22_X1 i_25_25_159 (.A1(\buffer[7][1][0] [15]), .A2(n_29), .B1(n_25), 
      .B2(\buffer[0][1][0] [15]), .ZN(n_25_25_143));
   AOI22_X1 i_25_25_160 (.A1(\buffer[15][1][0] [15]), .A2(n_22), .B1(n_27), 
      .B2(\buffer[12][1][0] [15]), .ZN(n_25_25_144));
   NAND4_X1 i_28_38_0 (.A1(n_28_38_8), .A2(n_28_38_6), .A3(n_28_38_4), .A4(
      n_28_38_0), .ZN(\output_filter[3][3] [0]));
   AOI221_X1 i_28_38_1 (.A(n_28_38_1), .B1(n_25), .B2(\buffer[0][3][3] [0]), 
      .C1(\buffer[12][3][3] [0]), .C2(n_27), .ZN(n_28_38_0));
   NAND4_X1 i_28_38_2 (.A1(n_28_38_7), .A2(n_28_38_5), .A3(n_28_38_3), .A4(
      n_28_38_2), .ZN(n_28_38_1));
   AOI22_X1 i_28_38_3 (.A1(\buffer[15][3][3] [0]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][3] [0]), .ZN(n_28_38_2));
   AOI22_X1 i_28_38_4 (.A1(\buffer[10][3][3] [0]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][3] [0]), .ZN(n_28_38_3));
   AOI22_X1 i_28_38_5 (.A1(\buffer[6][3][3] [0]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][3][3] [0]), .ZN(n_28_38_4));
   AOI22_X1 i_28_38_6 (.A1(\buffer[9][3][3] [0]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][3][3] [0]), .ZN(n_28_38_5));
   AOI22_X1 i_28_38_7 (.A1(\buffer[14][3][3] [0]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][3] [0]), .ZN(n_28_38_6));
   AOI22_X1 i_28_38_8 (.A1(\buffer[11][3][3] [0]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][3] [0]), .ZN(n_28_38_7));
   AOI22_X1 i_28_38_9 (.A1(\buffer[13][3][3] [0]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][3] [0]), .ZN(n_28_38_8));
   NAND4_X1 i_28_38_10 (.A1(n_28_38_17), .A2(n_28_38_15), .A3(n_28_38_13), 
      .A4(n_28_38_9), .ZN(\output_filter[3][3] [1]));
   AOI221_X1 i_28_38_11 (.A(n_28_38_10), .B1(n_25), .B2(\buffer[0][3][3] [1]), 
      .C1(\buffer[12][3][3] [1]), .C2(n_27), .ZN(n_28_38_9));
   NAND4_X1 i_28_38_12 (.A1(n_28_38_16), .A2(n_28_38_14), .A3(n_28_38_12), 
      .A4(n_28_38_11), .ZN(n_28_38_10));
   AOI22_X1 i_28_38_13 (.A1(\buffer[15][3][3] [1]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][3] [1]), .ZN(n_28_38_11));
   AOI22_X1 i_28_38_14 (.A1(\buffer[10][3][3] [1]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][3] [1]), .ZN(n_28_38_12));
   AOI22_X1 i_28_38_15 (.A1(\buffer[6][3][3] [1]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][3] [1]), .ZN(n_28_38_13));
   AOI22_X1 i_28_38_16 (.A1(\buffer[9][3][3] [1]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][3][3] [1]), .ZN(n_28_38_14));
   AOI22_X1 i_28_38_17 (.A1(\buffer[14][3][3] [1]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][3] [1]), .ZN(n_28_38_15));
   AOI22_X1 i_28_38_18 (.A1(\buffer[11][3][3] [1]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][3] [1]), .ZN(n_28_38_16));
   AOI22_X1 i_28_38_19 (.A1(\buffer[13][3][3] [1]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][3] [1]), .ZN(n_28_38_17));
   NAND4_X1 i_28_38_20 (.A1(n_28_38_26), .A2(n_28_38_24), .A3(n_28_38_22), 
      .A4(n_28_38_18), .ZN(\output_filter[3][3] [2]));
   AOI221_X1 i_28_38_21 (.A(n_28_38_19), .B1(n_25), .B2(\buffer[0][3][3] [2]), 
      .C1(\buffer[12][3][3] [2]), .C2(n_27), .ZN(n_28_38_18));
   NAND4_X1 i_28_38_22 (.A1(n_28_38_25), .A2(n_28_38_23), .A3(n_28_38_21), 
      .A4(n_28_38_20), .ZN(n_28_38_19));
   AOI22_X1 i_28_38_23 (.A1(\buffer[15][3][3] [2]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][3] [2]), .ZN(n_28_38_20));
   AOI22_X1 i_28_38_24 (.A1(\buffer[10][3][3] [2]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][3] [2]), .ZN(n_28_38_21));
   AOI22_X1 i_28_38_25 (.A1(\buffer[6][3][3] [2]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][3] [2]), .ZN(n_28_38_22));
   AOI22_X1 i_28_38_26 (.A1(\buffer[9][3][3] [2]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][3][3] [2]), .ZN(n_28_38_23));
   AOI22_X1 i_28_38_27 (.A1(\buffer[14][3][3] [2]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][3] [2]), .ZN(n_28_38_24));
   AOI22_X1 i_28_38_28 (.A1(\buffer[11][3][3] [2]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][3] [2]), .ZN(n_28_38_25));
   AOI22_X1 i_28_38_29 (.A1(\buffer[13][3][3] [2]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][3] [2]), .ZN(n_28_38_26));
   NAND4_X1 i_28_38_30 (.A1(n_28_38_35), .A2(n_28_38_33), .A3(n_28_38_31), 
      .A4(n_28_38_27), .ZN(\output_filter[3][3] [3]));
   AOI221_X1 i_28_38_31 (.A(n_28_38_28), .B1(n_25), .B2(\buffer[0][3][3] [3]), 
      .C1(\buffer[12][3][3] [3]), .C2(n_27), .ZN(n_28_38_27));
   NAND4_X1 i_28_38_32 (.A1(n_28_38_34), .A2(n_28_38_32), .A3(n_28_38_30), 
      .A4(n_28_38_29), .ZN(n_28_38_28));
   AOI22_X1 i_28_38_33 (.A1(\buffer[15][3][3] [3]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][3] [3]), .ZN(n_28_38_29));
   AOI22_X1 i_28_38_34 (.A1(\buffer[10][3][3] [3]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][3] [3]), .ZN(n_28_38_30));
   AOI22_X1 i_28_38_35 (.A1(\buffer[6][3][3] [3]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][3] [3]), .ZN(n_28_38_31));
   AOI22_X1 i_28_38_36 (.A1(\buffer[9][3][3] [3]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][3][3] [3]), .ZN(n_28_38_32));
   AOI22_X1 i_28_38_37 (.A1(\buffer[14][3][3] [3]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][3] [3]), .ZN(n_28_38_33));
   AOI22_X1 i_28_38_38 (.A1(\buffer[11][3][3] [3]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][3] [3]), .ZN(n_28_38_34));
   AOI22_X1 i_28_38_39 (.A1(\buffer[13][3][3] [3]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][3] [3]), .ZN(n_28_38_35));
   NAND4_X1 i_28_38_40 (.A1(n_28_38_44), .A2(n_28_38_42), .A3(n_28_38_40), 
      .A4(n_28_38_36), .ZN(\output_filter[3][3] [4]));
   AOI221_X1 i_28_38_41 (.A(n_28_38_37), .B1(n_25), .B2(\buffer[0][3][3] [4]), 
      .C1(\buffer[12][3][3] [4]), .C2(n_27), .ZN(n_28_38_36));
   NAND4_X1 i_28_38_42 (.A1(n_28_38_43), .A2(n_28_38_41), .A3(n_28_38_39), 
      .A4(n_28_38_38), .ZN(n_28_38_37));
   AOI22_X1 i_28_38_43 (.A1(\buffer[15][3][3] [4]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][3] [4]), .ZN(n_28_38_38));
   AOI22_X1 i_28_38_44 (.A1(\buffer[10][3][3] [4]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][3] [4]), .ZN(n_28_38_39));
   AOI22_X1 i_28_38_45 (.A1(\buffer[6][3][3] [4]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][3] [4]), .ZN(n_28_38_40));
   AOI22_X1 i_28_38_46 (.A1(\buffer[9][3][3] [4]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][3][3] [4]), .ZN(n_28_38_41));
   AOI22_X1 i_28_38_47 (.A1(\buffer[14][3][3] [4]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][3] [4]), .ZN(n_28_38_42));
   AOI22_X1 i_28_38_48 (.A1(\buffer[11][3][3] [4]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][3] [4]), .ZN(n_28_38_43));
   AOI22_X1 i_28_38_49 (.A1(\buffer[13][3][3] [4]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][3][3] [4]), .ZN(n_28_38_44));
   NAND4_X1 i_28_38_50 (.A1(n_28_38_53), .A2(n_28_38_51), .A3(n_28_38_49), 
      .A4(n_28_38_45), .ZN(\output_filter[3][3] [5]));
   AOI221_X1 i_28_38_51 (.A(n_28_38_46), .B1(n_25), .B2(\buffer[0][3][3] [5]), 
      .C1(\buffer[12][3][3] [5]), .C2(n_27), .ZN(n_28_38_45));
   NAND4_X1 i_28_38_52 (.A1(n_28_38_52), .A2(n_28_38_50), .A3(n_28_38_48), 
      .A4(n_28_38_47), .ZN(n_28_38_46));
   AOI22_X1 i_28_38_53 (.A1(\buffer[15][3][3] [5]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][3] [5]), .ZN(n_28_38_47));
   AOI22_X1 i_28_38_54 (.A1(\buffer[10][3][3] [5]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][3] [5]), .ZN(n_28_38_48));
   AOI22_X1 i_28_38_55 (.A1(\buffer[6][3][3] [5]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][3] [5]), .ZN(n_28_38_49));
   AOI22_X1 i_28_38_56 (.A1(\buffer[9][3][3] [5]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][3][3] [5]), .ZN(n_28_38_50));
   AOI22_X1 i_28_38_57 (.A1(\buffer[14][3][3] [5]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][3] [5]), .ZN(n_28_38_51));
   AOI22_X1 i_28_38_58 (.A1(\buffer[11][3][3] [5]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][3] [5]), .ZN(n_28_38_52));
   AOI22_X1 i_28_38_59 (.A1(\buffer[13][3][3] [5]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][3] [5]), .ZN(n_28_38_53));
   NAND4_X1 i_28_38_60 (.A1(n_28_38_62), .A2(n_28_38_60), .A3(n_28_38_58), 
      .A4(n_28_38_54), .ZN(\output_filter[3][3] [6]));
   AOI221_X1 i_28_38_61 (.A(n_28_38_55), .B1(n_25), .B2(\buffer[0][3][3] [6]), 
      .C1(\buffer[12][3][3] [6]), .C2(n_27), .ZN(n_28_38_54));
   NAND4_X1 i_28_38_62 (.A1(n_28_38_61), .A2(n_28_38_59), .A3(n_28_38_57), 
      .A4(n_28_38_56), .ZN(n_28_38_55));
   AOI22_X1 i_28_38_63 (.A1(\buffer[15][3][3] [6]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][3] [6]), .ZN(n_28_38_56));
   AOI22_X1 i_28_38_64 (.A1(\buffer[10][3][3] [6]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][3] [6]), .ZN(n_28_38_57));
   AOI22_X1 i_28_38_65 (.A1(\buffer[6][3][3] [6]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][3] [6]), .ZN(n_28_38_58));
   AOI22_X1 i_28_38_66 (.A1(\buffer[9][3][3] [6]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][3][3] [6]), .ZN(n_28_38_59));
   AOI22_X1 i_28_38_67 (.A1(\buffer[14][3][3] [6]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][3] [6]), .ZN(n_28_38_60));
   AOI22_X1 i_28_38_68 (.A1(\buffer[11][3][3] [6]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][3] [6]), .ZN(n_28_38_61));
   AOI22_X1 i_28_38_69 (.A1(\buffer[13][3][3] [6]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][3] [6]), .ZN(n_28_38_62));
   NAND4_X1 i_28_38_70 (.A1(n_28_38_71), .A2(n_28_38_69), .A3(n_28_38_67), 
      .A4(n_28_38_63), .ZN(\output_filter[3][3] [7]));
   AOI221_X1 i_28_38_71 (.A(n_28_38_64), .B1(n_25), .B2(\buffer[0][3][3] [7]), 
      .C1(\buffer[12][3][3] [7]), .C2(n_27), .ZN(n_28_38_63));
   NAND4_X1 i_28_38_72 (.A1(n_28_38_70), .A2(n_28_38_68), .A3(n_28_38_66), 
      .A4(n_28_38_65), .ZN(n_28_38_64));
   AOI22_X1 i_28_38_73 (.A1(\buffer[15][3][3] [7]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][3] [7]), .ZN(n_28_38_65));
   AOI22_X1 i_28_38_74 (.A1(\buffer[10][3][3] [7]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][3] [7]), .ZN(n_28_38_66));
   AOI22_X1 i_28_38_75 (.A1(\buffer[6][3][3] [7]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][3] [7]), .ZN(n_28_38_67));
   AOI22_X1 i_28_38_76 (.A1(\buffer[9][3][3] [7]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][3][3] [7]), .ZN(n_28_38_68));
   AOI22_X1 i_28_38_77 (.A1(\buffer[14][3][3] [7]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][3] [7]), .ZN(n_28_38_69));
   AOI22_X1 i_28_38_78 (.A1(\buffer[11][3][3] [7]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][3] [7]), .ZN(n_28_38_70));
   AOI22_X1 i_28_38_79 (.A1(\buffer[13][3][3] [7]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][3][3] [7]), .ZN(n_28_38_71));
   NAND4_X1 i_28_38_80 (.A1(n_28_38_80), .A2(n_28_38_78), .A3(n_28_38_76), 
      .A4(n_28_38_72), .ZN(\output_filter[3][3] [8]));
   AOI221_X1 i_28_38_81 (.A(n_28_38_73), .B1(n_25), .B2(\buffer[0][3][3] [8]), 
      .C1(\buffer[12][3][3] [8]), .C2(n_27), .ZN(n_28_38_72));
   NAND4_X1 i_28_38_82 (.A1(n_28_38_79), .A2(n_28_38_77), .A3(n_28_38_75), 
      .A4(n_28_38_74), .ZN(n_28_38_73));
   AOI22_X1 i_28_38_83 (.A1(\buffer[15][3][3] [8]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][3] [8]), .ZN(n_28_38_74));
   AOI22_X1 i_28_38_84 (.A1(\buffer[10][3][3] [8]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][3] [8]), .ZN(n_28_38_75));
   AOI22_X1 i_28_38_85 (.A1(\buffer[6][3][3] [8]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][3] [8]), .ZN(n_28_38_76));
   AOI22_X1 i_28_38_86 (.A1(\buffer[9][3][3] [8]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][3][3] [8]), .ZN(n_28_38_77));
   AOI22_X1 i_28_38_87 (.A1(\buffer[14][3][3] [8]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][3] [8]), .ZN(n_28_38_78));
   AOI22_X1 i_28_38_88 (.A1(\buffer[11][3][3] [8]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][3] [8]), .ZN(n_28_38_79));
   AOI22_X1 i_28_38_89 (.A1(\buffer[13][3][3] [8]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][3] [8]), .ZN(n_28_38_80));
   NAND4_X1 i_28_38_90 (.A1(n_28_38_89), .A2(n_28_38_87), .A3(n_28_38_85), 
      .A4(n_28_38_81), .ZN(\output_filter[3][3] [9]));
   AOI221_X1 i_28_38_91 (.A(n_28_38_82), .B1(n_25), .B2(\buffer[0][3][3] [9]), 
      .C1(\buffer[12][3][3] [9]), .C2(n_27), .ZN(n_28_38_81));
   NAND4_X1 i_28_38_92 (.A1(n_28_38_88), .A2(n_28_38_86), .A3(n_28_38_84), 
      .A4(n_28_38_83), .ZN(n_28_38_82));
   AOI22_X1 i_28_38_93 (.A1(\buffer[15][3][3] [9]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][3] [9]), .ZN(n_28_38_83));
   AOI22_X1 i_28_38_94 (.A1(\buffer[10][3][3] [9]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][3] [9]), .ZN(n_28_38_84));
   AOI22_X1 i_28_38_95 (.A1(\buffer[6][3][3] [9]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][3] [9]), .ZN(n_28_38_85));
   AOI22_X1 i_28_38_96 (.A1(\buffer[9][3][3] [9]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][3][3] [9]), .ZN(n_28_38_86));
   AOI22_X1 i_28_38_97 (.A1(\buffer[14][3][3] [9]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][3] [9]), .ZN(n_28_38_87));
   AOI22_X1 i_28_38_98 (.A1(\buffer[11][3][3] [9]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][3] [9]), .ZN(n_28_38_88));
   AOI22_X1 i_28_38_99 (.A1(\buffer[13][3][3] [9]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][3][3] [9]), .ZN(n_28_38_89));
   NAND4_X1 i_28_38_100 (.A1(n_28_38_98), .A2(n_28_38_96), .A3(n_28_38_94), 
      .A4(n_28_38_90), .ZN(\output_filter[3][3] [10]));
   AOI221_X1 i_28_38_101 (.A(n_28_38_91), .B1(n_25), .B2(\buffer[0][3][3] [10]), 
      .C1(\buffer[12][3][3] [10]), .C2(n_27), .ZN(n_28_38_90));
   NAND4_X1 i_28_38_102 (.A1(n_28_38_97), .A2(n_28_38_95), .A3(n_28_38_93), 
      .A4(n_28_38_92), .ZN(n_28_38_91));
   AOI22_X1 i_28_38_103 (.A1(\buffer[15][3][3] [10]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][3] [10]), .ZN(n_28_38_92));
   AOI22_X1 i_28_38_104 (.A1(\buffer[10][3][3] [10]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][3] [10]), .ZN(n_28_38_93));
   AOI22_X1 i_28_38_105 (.A1(\buffer[6][3][3] [10]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][3] [10]), .ZN(n_28_38_94));
   AOI22_X1 i_28_38_106 (.A1(\buffer[9][3][3] [10]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][3][3] [10]), .ZN(n_28_38_95));
   AOI22_X1 i_28_38_107 (.A1(\buffer[14][3][3] [10]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][3] [10]), .ZN(n_28_38_96));
   AOI22_X1 i_28_38_108 (.A1(\buffer[11][3][3] [10]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][3] [10]), .ZN(n_28_38_97));
   AOI22_X1 i_28_38_109 (.A1(\buffer[13][3][3] [10]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][3] [10]), .ZN(n_28_38_98));
   NAND4_X1 i_28_38_110 (.A1(n_28_38_107), .A2(n_28_38_105), .A3(n_28_38_103), 
      .A4(n_28_38_99), .ZN(\output_filter[3][3] [11]));
   AOI221_X1 i_28_38_111 (.A(n_28_38_100), .B1(n_25), .B2(\buffer[0][3][3] [11]), 
      .C1(\buffer[12][3][3] [11]), .C2(n_27), .ZN(n_28_38_99));
   NAND4_X1 i_28_38_112 (.A1(n_28_38_106), .A2(n_28_38_104), .A3(n_28_38_102), 
      .A4(n_28_38_101), .ZN(n_28_38_100));
   AOI22_X1 i_28_38_113 (.A1(\buffer[15][3][3] [11]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][3] [11]), .ZN(n_28_38_101));
   AOI22_X1 i_28_38_114 (.A1(\buffer[10][3][3] [11]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][3] [11]), .ZN(n_28_38_102));
   AOI22_X1 i_28_38_115 (.A1(\buffer[6][3][3] [11]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][3] [11]), .ZN(n_28_38_103));
   AOI22_X1 i_28_38_116 (.A1(\buffer[9][3][3] [11]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][3][3] [11]), .ZN(n_28_38_104));
   AOI22_X1 i_28_38_117 (.A1(\buffer[14][3][3] [11]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][3] [11]), .ZN(n_28_38_105));
   AOI22_X1 i_28_38_118 (.A1(\buffer[11][3][3] [11]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][3] [11]), .ZN(n_28_38_106));
   AOI22_X1 i_28_38_119 (.A1(\buffer[13][3][3] [11]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][3][3] [11]), .ZN(n_28_38_107));
   NAND4_X1 i_28_38_120 (.A1(n_28_38_116), .A2(n_28_38_114), .A3(n_28_38_112), 
      .A4(n_28_38_108), .ZN(\output_filter[3][3] [12]));
   AOI221_X1 i_28_38_121 (.A(n_28_38_109), .B1(n_25), .B2(\buffer[0][3][3] [12]), 
      .C1(\buffer[12][3][3] [12]), .C2(n_27), .ZN(n_28_38_108));
   NAND4_X1 i_28_38_122 (.A1(n_28_38_115), .A2(n_28_38_113), .A3(n_28_38_111), 
      .A4(n_28_38_110), .ZN(n_28_38_109));
   AOI22_X1 i_28_38_123 (.A1(\buffer[15][3][3] [12]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][3] [12]), .ZN(n_28_38_110));
   AOI22_X1 i_28_38_124 (.A1(\buffer[10][3][3] [12]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][3] [12]), .ZN(n_28_38_111));
   AOI22_X1 i_28_38_125 (.A1(\buffer[6][3][3] [12]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][3] [12]), .ZN(n_28_38_112));
   AOI22_X1 i_28_38_126 (.A1(\buffer[9][3][3] [12]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][3][3] [12]), .ZN(n_28_38_113));
   AOI22_X1 i_28_38_127 (.A1(\buffer[14][3][3] [12]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][3] [12]), .ZN(n_28_38_114));
   AOI22_X1 i_28_38_128 (.A1(\buffer[11][3][3] [12]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][3] [12]), .ZN(n_28_38_115));
   AOI22_X1 i_28_38_129 (.A1(\buffer[13][3][3] [12]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][3] [12]), .ZN(n_28_38_116));
   NAND4_X1 i_28_38_130 (.A1(n_28_38_125), .A2(n_28_38_123), .A3(n_28_38_121), 
      .A4(n_28_38_117), .ZN(\output_filter[3][3] [13]));
   AOI221_X1 i_28_38_131 (.A(n_28_38_118), .B1(n_25), .B2(\buffer[0][3][3] [13]), 
      .C1(\buffer[12][3][3] [13]), .C2(n_27), .ZN(n_28_38_117));
   NAND4_X1 i_28_38_132 (.A1(n_28_38_124), .A2(n_28_38_122), .A3(n_28_38_120), 
      .A4(n_28_38_119), .ZN(n_28_38_118));
   AOI22_X1 i_28_38_133 (.A1(\buffer[15][3][3] [13]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][3][3] [13]), .ZN(n_28_38_119));
   AOI22_X1 i_28_38_134 (.A1(\buffer[10][3][3] [13]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][3][3] [13]), .ZN(n_28_38_120));
   AOI22_X1 i_28_38_135 (.A1(\buffer[6][3][3] [13]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][3] [13]), .ZN(n_28_38_121));
   AOI22_X1 i_28_38_136 (.A1(\buffer[9][3][3] [13]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][3][3] [13]), .ZN(n_28_38_122));
   AOI22_X1 i_28_38_137 (.A1(\buffer[14][3][3] [13]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][3] [13]), .ZN(n_28_38_123));
   AOI22_X1 i_28_38_138 (.A1(\buffer[11][3][3] [13]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][3] [13]), .ZN(n_28_38_124));
   AOI22_X1 i_28_38_139 (.A1(\buffer[13][3][3] [13]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][3][3] [13]), .ZN(n_28_38_125));
   NAND4_X1 i_28_38_140 (.A1(n_28_38_134), .A2(n_28_38_132), .A3(n_28_38_130), 
      .A4(n_28_38_126), .ZN(\output_filter[3][3] [14]));
   AOI221_X1 i_28_38_141 (.A(n_28_38_127), .B1(n_25), .B2(\buffer[0][3][3] [14]), 
      .C1(\buffer[12][3][3] [14]), .C2(n_27), .ZN(n_28_38_126));
   NAND4_X1 i_28_38_142 (.A1(n_28_38_133), .A2(n_28_38_131), .A3(n_28_38_129), 
      .A4(n_28_38_128), .ZN(n_28_38_127));
   AOI22_X1 i_28_38_143 (.A1(\buffer[15][3][3] [14]), .A2(n_22), .B1(n_16), 
      .B2(\buffer[8][3][3] [14]), .ZN(n_28_38_128));
   AOI22_X1 i_28_38_144 (.A1(\buffer[10][3][3] [14]), .A2(n_21), .B1(n_29), 
      .B2(\buffer[7][3][3] [14]), .ZN(n_28_38_129));
   AOI22_X1 i_28_38_145 (.A1(\buffer[6][3][3] [14]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][3][3] [14]), .ZN(n_28_38_130));
   AOI22_X1 i_28_38_146 (.A1(\buffer[9][3][3] [14]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][3][3] [14]), .ZN(n_28_38_131));
   AOI22_X1 i_28_38_147 (.A1(\buffer[14][3][3] [14]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][3][3] [14]), .ZN(n_28_38_132));
   AOI22_X1 i_28_38_148 (.A1(\buffer[11][3][3] [14]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][3][3] [14]), .ZN(n_28_38_133));
   AOI22_X1 i_28_38_149 (.A1(\buffer[13][3][3] [14]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][3][3] [14]), .ZN(n_28_38_134));
   NAND2_X1 i_28_38_150 (.A1(n_28_38_137), .A2(n_28_38_135), .ZN(
      \output_filter[3][3] [15]));
   AOI221_X1 i_28_38_151 (.A(n_28_38_136), .B1(n_31), .B2(\buffer[3][3][3] [15]), 
      .C1(\buffer[14][3][3] [15]), .C2(n_19), .ZN(n_28_38_135));
   NAND3_X1 i_28_38_152 (.A1(n_28_38_143), .A2(n_28_38_141), .A3(n_28_38_139), 
      .ZN(n_28_38_136));
   AOI221_X1 i_28_38_153 (.A(n_28_38_138), .B1(n_16), .B2(\buffer[8][3][3] [15]), 
      .C1(\buffer[13][3][3] [15]), .C2(n_26), .ZN(n_28_38_137));
   NAND3_X1 i_28_38_154 (.A1(n_28_38_144), .A2(n_28_38_142), .A3(n_28_38_140), 
      .ZN(n_28_38_138));
   AOI22_X1 i_28_38_155 (.A1(\buffer[11][3][3] [15]), .A2(n_17), .B1(n_24), 
      .B2(\buffer[2][3][3] [15]), .ZN(n_28_38_139));
   AOI22_X1 i_28_38_156 (.A1(\buffer[10][3][3] [15]), .A2(n_21), .B1(n_23), 
      .B2(\buffer[1][3][3] [15]), .ZN(n_28_38_140));
   AOI22_X1 i_28_38_157 (.A1(\buffer[6][3][3] [15]), .A2(n_28), .B1(n_18), 
      .B2(\buffer[5][3][3] [15]), .ZN(n_28_38_141));
   AOI22_X1 i_28_38_158 (.A1(\buffer[9][3][3] [15]), .A2(n_20), .B1(n_30), 
      .B2(\buffer[4][3][3] [15]), .ZN(n_28_38_142));
   AOI22_X1 i_28_38_159 (.A1(\buffer[7][3][3] [15]), .A2(n_29), .B1(n_25), 
      .B2(\buffer[0][3][3] [15]), .ZN(n_28_38_143));
   AOI22_X1 i_28_38_160 (.A1(\buffer[15][3][3] [15]), .A2(n_22), .B1(n_27), 
      .B2(\buffer[12][3][3] [15]), .ZN(n_28_38_144));
   NAND4_X1 i_24_24_0 (.A1(n_24_24_8), .A2(n_24_24_6), .A3(n_24_24_4), .A4(
      n_24_24_0), .ZN(\output_filter[0][4] [0]));
   AOI221_X1 i_24_24_1 (.A(n_24_24_1), .B1(n_25), .B2(\buffer[0][0][4] [0]), 
      .C1(\buffer[12][0][4] [0]), .C2(n_27), .ZN(n_24_24_0));
   NAND4_X1 i_24_24_2 (.A1(n_24_24_7), .A2(n_24_24_5), .A3(n_24_24_3), .A4(
      n_24_24_2), .ZN(n_24_24_1));
   AOI22_X1 i_24_24_3 (.A1(\buffer[15][0][4] [0]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][4] [0]), .ZN(n_24_24_2));
   AOI22_X1 i_24_24_4 (.A1(\buffer[10][0][4] [0]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][4] [0]), .ZN(n_24_24_3));
   AOI22_X1 i_24_24_5 (.A1(\buffer[6][0][4] [0]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][0][4] [0]), .ZN(n_24_24_4));
   AOI22_X1 i_24_24_6 (.A1(\buffer[9][0][4] [0]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][0][4] [0]), .ZN(n_24_24_5));
   AOI22_X1 i_24_24_7 (.A1(\buffer[14][0][4] [0]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][4] [0]), .ZN(n_24_24_6));
   AOI22_X1 i_24_24_8 (.A1(\buffer[11][0][4] [0]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][4] [0]), .ZN(n_24_24_7));
   AOI22_X1 i_24_24_9 (.A1(\buffer[13][0][4] [0]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][4] [0]), .ZN(n_24_24_8));
   NAND4_X1 i_24_24_10 (.A1(n_24_24_17), .A2(n_24_24_15), .A3(n_24_24_13), 
      .A4(n_24_24_9), .ZN(\output_filter[0][4] [1]));
   AOI221_X1 i_24_24_11 (.A(n_24_24_10), .B1(n_25), .B2(\buffer[0][0][4] [1]), 
      .C1(\buffer[12][0][4] [1]), .C2(n_27), .ZN(n_24_24_9));
   NAND4_X1 i_24_24_12 (.A1(n_24_24_16), .A2(n_24_24_14), .A3(n_24_24_12), 
      .A4(n_24_24_11), .ZN(n_24_24_10));
   AOI22_X1 i_24_24_13 (.A1(\buffer[15][0][4] [1]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][4] [1]), .ZN(n_24_24_11));
   AOI22_X1 i_24_24_14 (.A1(\buffer[10][0][4] [1]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][4] [1]), .ZN(n_24_24_12));
   AOI22_X1 i_24_24_15 (.A1(\buffer[6][0][4] [1]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][4] [1]), .ZN(n_24_24_13));
   AOI22_X1 i_24_24_16 (.A1(\buffer[9][0][4] [1]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][4] [1]), .ZN(n_24_24_14));
   AOI22_X1 i_24_24_17 (.A1(\buffer[14][0][4] [1]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][4] [1]), .ZN(n_24_24_15));
   AOI22_X1 i_24_24_18 (.A1(\buffer[11][0][4] [1]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][4] [1]), .ZN(n_24_24_16));
   AOI22_X1 i_24_24_19 (.A1(\buffer[13][0][4] [1]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][4] [1]), .ZN(n_24_24_17));
   NAND4_X1 i_24_24_20 (.A1(n_24_24_26), .A2(n_24_24_24), .A3(n_24_24_22), 
      .A4(n_24_24_18), .ZN(\output_filter[0][4] [2]));
   AOI221_X1 i_24_24_21 (.A(n_24_24_19), .B1(n_25), .B2(\buffer[0][0][4] [2]), 
      .C1(\buffer[12][0][4] [2]), .C2(n_27), .ZN(n_24_24_18));
   NAND4_X1 i_24_24_22 (.A1(n_24_24_25), .A2(n_24_24_23), .A3(n_24_24_21), 
      .A4(n_24_24_20), .ZN(n_24_24_19));
   AOI22_X1 i_24_24_23 (.A1(\buffer[15][0][4] [2]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][4] [2]), .ZN(n_24_24_20));
   AOI22_X1 i_24_24_24 (.A1(\buffer[10][0][4] [2]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][4] [2]), .ZN(n_24_24_21));
   AOI22_X1 i_24_24_25 (.A1(\buffer[6][0][4] [2]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][4] [2]), .ZN(n_24_24_22));
   AOI22_X1 i_24_24_26 (.A1(\buffer[9][0][4] [2]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][4] [2]), .ZN(n_24_24_23));
   AOI22_X1 i_24_24_27 (.A1(\buffer[14][0][4] [2]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][4] [2]), .ZN(n_24_24_24));
   AOI22_X1 i_24_24_28 (.A1(\buffer[11][0][4] [2]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][4] [2]), .ZN(n_24_24_25));
   AOI22_X1 i_24_24_29 (.A1(\buffer[13][0][4] [2]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][4] [2]), .ZN(n_24_24_26));
   NAND4_X1 i_24_24_30 (.A1(n_24_24_35), .A2(n_24_24_33), .A3(n_24_24_31), 
      .A4(n_24_24_27), .ZN(\output_filter[0][4] [3]));
   AOI221_X1 i_24_24_31 (.A(n_24_24_28), .B1(n_25), .B2(\buffer[0][0][4] [3]), 
      .C1(\buffer[12][0][4] [3]), .C2(n_27), .ZN(n_24_24_27));
   NAND4_X1 i_24_24_32 (.A1(n_24_24_34), .A2(n_24_24_32), .A3(n_24_24_30), 
      .A4(n_24_24_29), .ZN(n_24_24_28));
   AOI22_X1 i_24_24_33 (.A1(\buffer[15][0][4] [3]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][4] [3]), .ZN(n_24_24_29));
   AOI22_X1 i_24_24_34 (.A1(\buffer[10][0][4] [3]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][4] [3]), .ZN(n_24_24_30));
   AOI22_X1 i_24_24_35 (.A1(\buffer[6][0][4] [3]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][4] [3]), .ZN(n_24_24_31));
   AOI22_X1 i_24_24_36 (.A1(\buffer[9][0][4] [3]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][4] [3]), .ZN(n_24_24_32));
   AOI22_X1 i_24_24_37 (.A1(\buffer[14][0][4] [3]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][4] [3]), .ZN(n_24_24_33));
   AOI22_X1 i_24_24_38 (.A1(\buffer[11][0][4] [3]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][4] [3]), .ZN(n_24_24_34));
   AOI22_X1 i_24_24_39 (.A1(\buffer[13][0][4] [3]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][4] [3]), .ZN(n_24_24_35));
   NAND4_X1 i_24_24_40 (.A1(n_24_24_44), .A2(n_24_24_42), .A3(n_24_24_40), 
      .A4(n_24_24_36), .ZN(\output_filter[0][4] [4]));
   AOI221_X1 i_24_24_41 (.A(n_24_24_37), .B1(n_25), .B2(\buffer[0][0][4] [4]), 
      .C1(\buffer[12][0][4] [4]), .C2(n_27), .ZN(n_24_24_36));
   NAND4_X1 i_24_24_42 (.A1(n_24_24_43), .A2(n_24_24_41), .A3(n_24_24_39), 
      .A4(n_24_24_38), .ZN(n_24_24_37));
   AOI22_X1 i_24_24_43 (.A1(\buffer[15][0][4] [4]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][4] [4]), .ZN(n_24_24_38));
   AOI22_X1 i_24_24_44 (.A1(\buffer[10][0][4] [4]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][4] [4]), .ZN(n_24_24_39));
   AOI22_X1 i_24_24_45 (.A1(\buffer[6][0][4] [4]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][4] [4]), .ZN(n_24_24_40));
   AOI22_X1 i_24_24_46 (.A1(\buffer[9][0][4] [4]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][0][4] [4]), .ZN(n_24_24_41));
   AOI22_X1 i_24_24_47 (.A1(\buffer[14][0][4] [4]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][4] [4]), .ZN(n_24_24_42));
   AOI22_X1 i_24_24_48 (.A1(\buffer[11][0][4] [4]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][4] [4]), .ZN(n_24_24_43));
   AOI22_X1 i_24_24_49 (.A1(\buffer[13][0][4] [4]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][0][4] [4]), .ZN(n_24_24_44));
   NAND4_X1 i_24_24_50 (.A1(n_24_24_53), .A2(n_24_24_51), .A3(n_24_24_49), 
      .A4(n_24_24_45), .ZN(\output_filter[0][4] [5]));
   AOI221_X1 i_24_24_51 (.A(n_24_24_46), .B1(n_25), .B2(\buffer[0][0][4] [5]), 
      .C1(\buffer[12][0][4] [5]), .C2(n_27), .ZN(n_24_24_45));
   NAND4_X1 i_24_24_52 (.A1(n_24_24_52), .A2(n_24_24_50), .A3(n_24_24_48), 
      .A4(n_24_24_47), .ZN(n_24_24_46));
   AOI22_X1 i_24_24_53 (.A1(\buffer[15][0][4] [5]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][4] [5]), .ZN(n_24_24_47));
   AOI22_X1 i_24_24_54 (.A1(\buffer[10][0][4] [5]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][4] [5]), .ZN(n_24_24_48));
   AOI22_X1 i_24_24_55 (.A1(\buffer[6][0][4] [5]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][4] [5]), .ZN(n_24_24_49));
   AOI22_X1 i_24_24_56 (.A1(\buffer[9][0][4] [5]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][4] [5]), .ZN(n_24_24_50));
   AOI22_X1 i_24_24_57 (.A1(\buffer[14][0][4] [5]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][4] [5]), .ZN(n_24_24_51));
   AOI22_X1 i_24_24_58 (.A1(\buffer[11][0][4] [5]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][4] [5]), .ZN(n_24_24_52));
   AOI22_X1 i_24_24_59 (.A1(\buffer[13][0][4] [5]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][4] [5]), .ZN(n_24_24_53));
   NAND4_X1 i_24_24_60 (.A1(n_24_24_62), .A2(n_24_24_60), .A3(n_24_24_58), 
      .A4(n_24_24_54), .ZN(\output_filter[0][4] [6]));
   AOI221_X1 i_24_24_61 (.A(n_24_24_55), .B1(n_25), .B2(\buffer[0][0][4] [6]), 
      .C1(\buffer[12][0][4] [6]), .C2(n_27), .ZN(n_24_24_54));
   NAND4_X1 i_24_24_62 (.A1(n_24_24_61), .A2(n_24_24_59), .A3(n_24_24_57), 
      .A4(n_24_24_56), .ZN(n_24_24_55));
   AOI22_X1 i_24_24_63 (.A1(\buffer[15][0][4] [6]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][4] [6]), .ZN(n_24_24_56));
   AOI22_X1 i_24_24_64 (.A1(\buffer[10][0][4] [6]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][4] [6]), .ZN(n_24_24_57));
   AOI22_X1 i_24_24_65 (.A1(\buffer[6][0][4] [6]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][4] [6]), .ZN(n_24_24_58));
   AOI22_X1 i_24_24_66 (.A1(\buffer[9][0][4] [6]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][4] [6]), .ZN(n_24_24_59));
   AOI22_X1 i_24_24_67 (.A1(\buffer[14][0][4] [6]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][4] [6]), .ZN(n_24_24_60));
   AOI22_X1 i_24_24_68 (.A1(\buffer[11][0][4] [6]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][4] [6]), .ZN(n_24_24_61));
   AOI22_X1 i_24_24_69 (.A1(\buffer[13][0][4] [6]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][4] [6]), .ZN(n_24_24_62));
   NAND4_X1 i_24_24_70 (.A1(n_24_24_71), .A2(n_24_24_69), .A3(n_24_24_67), 
      .A4(n_24_24_63), .ZN(\output_filter[0][4] [7]));
   AOI221_X1 i_24_24_71 (.A(n_24_24_64), .B1(n_25), .B2(\buffer[0][0][4] [7]), 
      .C1(\buffer[12][0][4] [7]), .C2(n_27), .ZN(n_24_24_63));
   NAND4_X1 i_24_24_72 (.A1(n_24_24_70), .A2(n_24_24_68), .A3(n_24_24_66), 
      .A4(n_24_24_65), .ZN(n_24_24_64));
   AOI22_X1 i_24_24_73 (.A1(\buffer[15][0][4] [7]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][4] [7]), .ZN(n_24_24_65));
   AOI22_X1 i_24_24_74 (.A1(\buffer[10][0][4] [7]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][4] [7]), .ZN(n_24_24_66));
   AOI22_X1 i_24_24_75 (.A1(\buffer[6][0][4] [7]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][4] [7]), .ZN(n_24_24_67));
   AOI22_X1 i_24_24_76 (.A1(\buffer[9][0][4] [7]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][0][4] [7]), .ZN(n_24_24_68));
   AOI22_X1 i_24_24_77 (.A1(\buffer[14][0][4] [7]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][4] [7]), .ZN(n_24_24_69));
   AOI22_X1 i_24_24_78 (.A1(\buffer[11][0][4] [7]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][4] [7]), .ZN(n_24_24_70));
   AOI22_X1 i_24_24_79 (.A1(\buffer[13][0][4] [7]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][0][4] [7]), .ZN(n_24_24_71));
   NAND4_X1 i_24_24_80 (.A1(n_24_24_80), .A2(n_24_24_78), .A3(n_24_24_76), 
      .A4(n_24_24_72), .ZN(\output_filter[0][4] [8]));
   AOI221_X1 i_24_24_81 (.A(n_24_24_73), .B1(n_25), .B2(\buffer[0][0][4] [8]), 
      .C1(\buffer[12][0][4] [8]), .C2(n_27), .ZN(n_24_24_72));
   NAND4_X1 i_24_24_82 (.A1(n_24_24_79), .A2(n_24_24_77), .A3(n_24_24_75), 
      .A4(n_24_24_74), .ZN(n_24_24_73));
   AOI22_X1 i_24_24_83 (.A1(\buffer[15][0][4] [8]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][4] [8]), .ZN(n_24_24_74));
   AOI22_X1 i_24_24_84 (.A1(\buffer[10][0][4] [8]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][4] [8]), .ZN(n_24_24_75));
   AOI22_X1 i_24_24_85 (.A1(\buffer[6][0][4] [8]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][4] [8]), .ZN(n_24_24_76));
   AOI22_X1 i_24_24_86 (.A1(\buffer[9][0][4] [8]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][4] [8]), .ZN(n_24_24_77));
   AOI22_X1 i_24_24_87 (.A1(\buffer[14][0][4] [8]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][4] [8]), .ZN(n_24_24_78));
   AOI22_X1 i_24_24_88 (.A1(\buffer[11][0][4] [8]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][4] [8]), .ZN(n_24_24_79));
   AOI22_X1 i_24_24_89 (.A1(\buffer[13][0][4] [8]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][4] [8]), .ZN(n_24_24_80));
   NAND4_X1 i_24_24_90 (.A1(n_24_24_89), .A2(n_24_24_87), .A3(n_24_24_85), 
      .A4(n_24_24_81), .ZN(\output_filter[0][4] [9]));
   AOI221_X1 i_24_24_91 (.A(n_24_24_82), .B1(n_25), .B2(\buffer[0][0][4] [9]), 
      .C1(\buffer[12][0][4] [9]), .C2(n_27), .ZN(n_24_24_81));
   NAND4_X1 i_24_24_92 (.A1(n_24_24_88), .A2(n_24_24_86), .A3(n_24_24_84), 
      .A4(n_24_24_83), .ZN(n_24_24_82));
   AOI22_X1 i_24_24_93 (.A1(\buffer[15][0][4] [9]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][4] [9]), .ZN(n_24_24_83));
   AOI22_X1 i_24_24_94 (.A1(\buffer[10][0][4] [9]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][4] [9]), .ZN(n_24_24_84));
   AOI22_X1 i_24_24_95 (.A1(\buffer[6][0][4] [9]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][4] [9]), .ZN(n_24_24_85));
   AOI22_X1 i_24_24_96 (.A1(\buffer[9][0][4] [9]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][0][4] [9]), .ZN(n_24_24_86));
   AOI22_X1 i_24_24_97 (.A1(\buffer[14][0][4] [9]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][4] [9]), .ZN(n_24_24_87));
   AOI22_X1 i_24_24_98 (.A1(\buffer[11][0][4] [9]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][4] [9]), .ZN(n_24_24_88));
   AOI22_X1 i_24_24_99 (.A1(\buffer[13][0][4] [9]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][0][4] [9]), .ZN(n_24_24_89));
   NAND4_X1 i_24_24_100 (.A1(n_24_24_98), .A2(n_24_24_96), .A3(n_24_24_94), 
      .A4(n_24_24_90), .ZN(\output_filter[0][4] [10]));
   AOI221_X1 i_24_24_101 (.A(n_24_24_91), .B1(n_25), .B2(\buffer[0][0][4] [10]), 
      .C1(\buffer[12][0][4] [10]), .C2(n_27), .ZN(n_24_24_90));
   NAND4_X1 i_24_24_102 (.A1(n_24_24_97), .A2(n_24_24_95), .A3(n_24_24_93), 
      .A4(n_24_24_92), .ZN(n_24_24_91));
   AOI22_X1 i_24_24_103 (.A1(\buffer[15][0][4] [10]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][4] [10]), .ZN(n_24_24_92));
   AOI22_X1 i_24_24_104 (.A1(\buffer[10][0][4] [10]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][4] [10]), .ZN(n_24_24_93));
   AOI22_X1 i_24_24_105 (.A1(\buffer[6][0][4] [10]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][4] [10]), .ZN(n_24_24_94));
   AOI22_X1 i_24_24_106 (.A1(\buffer[9][0][4] [10]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][4] [10]), .ZN(n_24_24_95));
   AOI22_X1 i_24_24_107 (.A1(\buffer[14][0][4] [10]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][4] [10]), .ZN(n_24_24_96));
   AOI22_X1 i_24_24_108 (.A1(\buffer[11][0][4] [10]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][4] [10]), .ZN(n_24_24_97));
   AOI22_X1 i_24_24_109 (.A1(\buffer[13][0][4] [10]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][4] [10]), .ZN(n_24_24_98));
   NAND4_X1 i_24_24_110 (.A1(n_24_24_107), .A2(n_24_24_105), .A3(n_24_24_103), 
      .A4(n_24_24_99), .ZN(\output_filter[0][4] [11]));
   AOI221_X1 i_24_24_111 (.A(n_24_24_100), .B1(n_25), .B2(\buffer[0][0][4] [11]), 
      .C1(\buffer[12][0][4] [11]), .C2(n_27), .ZN(n_24_24_99));
   NAND4_X1 i_24_24_112 (.A1(n_24_24_106), .A2(n_24_24_104), .A3(n_24_24_102), 
      .A4(n_24_24_101), .ZN(n_24_24_100));
   AOI22_X1 i_24_24_113 (.A1(\buffer[15][0][4] [11]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][4] [11]), .ZN(n_24_24_101));
   AOI22_X1 i_24_24_114 (.A1(\buffer[10][0][4] [11]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][4] [11]), .ZN(n_24_24_102));
   AOI22_X1 i_24_24_115 (.A1(\buffer[6][0][4] [11]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][4] [11]), .ZN(n_24_24_103));
   AOI22_X1 i_24_24_116 (.A1(\buffer[9][0][4] [11]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][0][4] [11]), .ZN(n_24_24_104));
   AOI22_X1 i_24_24_117 (.A1(\buffer[14][0][4] [11]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][4] [11]), .ZN(n_24_24_105));
   AOI22_X1 i_24_24_118 (.A1(\buffer[11][0][4] [11]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][4] [11]), .ZN(n_24_24_106));
   AOI22_X1 i_24_24_119 (.A1(\buffer[13][0][4] [11]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][0][4] [11]), .ZN(n_24_24_107));
   NAND4_X1 i_24_24_120 (.A1(n_24_24_116), .A2(n_24_24_114), .A3(n_24_24_112), 
      .A4(n_24_24_108), .ZN(\output_filter[0][4] [12]));
   AOI221_X1 i_24_24_121 (.A(n_24_24_109), .B1(n_25), .B2(\buffer[0][0][4] [12]), 
      .C1(\buffer[12][0][4] [12]), .C2(n_27), .ZN(n_24_24_108));
   NAND4_X1 i_24_24_122 (.A1(n_24_24_115), .A2(n_24_24_113), .A3(n_24_24_111), 
      .A4(n_24_24_110), .ZN(n_24_24_109));
   AOI22_X1 i_24_24_123 (.A1(\buffer[15][0][4] [12]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][4] [12]), .ZN(n_24_24_110));
   AOI22_X1 i_24_24_124 (.A1(\buffer[10][0][4] [12]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][4] [12]), .ZN(n_24_24_111));
   AOI22_X1 i_24_24_125 (.A1(\buffer[6][0][4] [12]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][4] [12]), .ZN(n_24_24_112));
   AOI22_X1 i_24_24_126 (.A1(\buffer[9][0][4] [12]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][4] [12]), .ZN(n_24_24_113));
   AOI22_X1 i_24_24_127 (.A1(\buffer[14][0][4] [12]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][4] [12]), .ZN(n_24_24_114));
   AOI22_X1 i_24_24_128 (.A1(\buffer[11][0][4] [12]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][4] [12]), .ZN(n_24_24_115));
   AOI22_X1 i_24_24_129 (.A1(\buffer[13][0][4] [12]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][4] [12]), .ZN(n_24_24_116));
   NAND4_X1 i_24_24_130 (.A1(n_24_24_125), .A2(n_24_24_123), .A3(n_24_24_121), 
      .A4(n_24_24_117), .ZN(\output_filter[0][4] [13]));
   AOI221_X1 i_24_24_131 (.A(n_24_24_118), .B1(n_25), .B2(\buffer[0][0][4] [13]), 
      .C1(\buffer[12][0][4] [13]), .C2(n_27), .ZN(n_24_24_117));
   NAND4_X1 i_24_24_132 (.A1(n_24_24_124), .A2(n_24_24_122), .A3(n_24_24_120), 
      .A4(n_24_24_119), .ZN(n_24_24_118));
   AOI22_X1 i_24_24_133 (.A1(\buffer[15][0][4] [13]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][4] [13]), .ZN(n_24_24_119));
   AOI22_X1 i_24_24_134 (.A1(\buffer[10][0][4] [13]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][4] [13]), .ZN(n_24_24_120));
   AOI22_X1 i_24_24_135 (.A1(\buffer[6][0][4] [13]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][4] [13]), .ZN(n_24_24_121));
   AOI22_X1 i_24_24_136 (.A1(\buffer[9][0][4] [13]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][0][4] [13]), .ZN(n_24_24_122));
   AOI22_X1 i_24_24_137 (.A1(\buffer[14][0][4] [13]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][4] [13]), .ZN(n_24_24_123));
   AOI22_X1 i_24_24_138 (.A1(\buffer[11][0][4] [13]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][4] [13]), .ZN(n_24_24_124));
   AOI22_X1 i_24_24_139 (.A1(\buffer[13][0][4] [13]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][0][4] [13]), .ZN(n_24_24_125));
   NAND4_X1 i_24_24_140 (.A1(n_24_24_134), .A2(n_24_24_132), .A3(n_24_24_130), 
      .A4(n_24_24_126), .ZN(\output_filter[0][4] [14]));
   AOI221_X1 i_24_24_141 (.A(n_24_24_127), .B1(n_25), .B2(\buffer[0][0][4] [14]), 
      .C1(\buffer[12][0][4] [14]), .C2(n_27), .ZN(n_24_24_126));
   NAND4_X1 i_24_24_142 (.A1(n_24_24_133), .A2(n_24_24_131), .A3(n_24_24_129), 
      .A4(n_24_24_128), .ZN(n_24_24_127));
   AOI22_X1 i_24_24_143 (.A1(\buffer[15][0][4] [14]), .A2(n_22), .B1(n_16), 
      .B2(\buffer[8][0][4] [14]), .ZN(n_24_24_128));
   AOI22_X1 i_24_24_144 (.A1(\buffer[10][0][4] [14]), .A2(n_21), .B1(n_29), 
      .B2(\buffer[7][0][4] [14]), .ZN(n_24_24_129));
   AOI22_X1 i_24_24_145 (.A1(\buffer[6][0][4] [14]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][4] [14]), .ZN(n_24_24_130));
   AOI22_X1 i_24_24_146 (.A1(\buffer[9][0][4] [14]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][4] [14]), .ZN(n_24_24_131));
   AOI22_X1 i_24_24_147 (.A1(\buffer[14][0][4] [14]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][4] [14]), .ZN(n_24_24_132));
   AOI22_X1 i_24_24_148 (.A1(\buffer[11][0][4] [14]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][4] [14]), .ZN(n_24_24_133));
   AOI22_X1 i_24_24_149 (.A1(\buffer[13][0][4] [14]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][4] [14]), .ZN(n_24_24_134));
   NAND2_X1 i_24_24_150 (.A1(n_24_24_137), .A2(n_24_24_135), .ZN(
      \output_filter[0][4] [15]));
   AOI221_X1 i_24_24_151 (.A(n_24_24_136), .B1(n_31), .B2(\buffer[3][0][4] [15]), 
      .C1(\buffer[14][0][4] [15]), .C2(n_19), .ZN(n_24_24_135));
   NAND3_X1 i_24_24_152 (.A1(n_24_24_143), .A2(n_24_24_141), .A3(n_24_24_139), 
      .ZN(n_24_24_136));
   AOI221_X1 i_24_24_153 (.A(n_24_24_138), .B1(n_16), .B2(\buffer[8][0][4] [15]), 
      .C1(\buffer[13][0][4] [15]), .C2(n_26), .ZN(n_24_24_137));
   NAND3_X1 i_24_24_154 (.A1(n_24_24_144), .A2(n_24_24_142), .A3(n_24_24_140), 
      .ZN(n_24_24_138));
   AOI22_X1 i_24_24_155 (.A1(\buffer[11][0][4] [15]), .A2(n_17), .B1(n_24), 
      .B2(\buffer[2][0][4] [15]), .ZN(n_24_24_139));
   AOI22_X1 i_24_24_156 (.A1(\buffer[10][0][4] [15]), .A2(n_21), .B1(n_23), 
      .B2(\buffer[1][0][4] [15]), .ZN(n_24_24_140));
   AOI22_X1 i_24_24_157 (.A1(\buffer[6][0][4] [15]), .A2(n_28), .B1(n_18), 
      .B2(\buffer[5][0][4] [15]), .ZN(n_24_24_141));
   AOI22_X1 i_24_24_158 (.A1(\buffer[9][0][4] [15]), .A2(n_20), .B1(n_30), 
      .B2(\buffer[4][0][4] [15]), .ZN(n_24_24_142));
   AOI22_X1 i_24_24_159 (.A1(\buffer[7][0][4] [15]), .A2(n_29), .B1(n_25), 
      .B2(\buffer[0][0][4] [15]), .ZN(n_24_24_143));
   AOI22_X1 i_24_24_160 (.A1(\buffer[15][0][4] [15]), .A2(n_22), .B1(n_27), 
      .B2(\buffer[12][0][4] [15]), .ZN(n_24_24_144));
   NAND4_X1 i_23_23_0 (.A1(n_23_23_8), .A2(n_23_23_6), .A3(n_23_23_4), .A4(
      n_23_23_0), .ZN(\output_filter[0][3] [0]));
   AOI221_X1 i_23_23_1 (.A(n_23_23_1), .B1(n_25), .B2(\buffer[0][0][3] [0]), 
      .C1(\buffer[12][0][3] [0]), .C2(n_27), .ZN(n_23_23_0));
   NAND4_X1 i_23_23_2 (.A1(n_23_23_7), .A2(n_23_23_5), .A3(n_23_23_3), .A4(
      n_23_23_2), .ZN(n_23_23_1));
   AOI22_X1 i_23_23_3 (.A1(\buffer[15][0][3] [0]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][3] [0]), .ZN(n_23_23_2));
   AOI22_X1 i_23_23_4 (.A1(\buffer[10][0][3] [0]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][3] [0]), .ZN(n_23_23_3));
   AOI22_X1 i_23_23_5 (.A1(\buffer[6][0][3] [0]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][0][3] [0]), .ZN(n_23_23_4));
   AOI22_X1 i_23_23_6 (.A1(\buffer[9][0][3] [0]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][0][3] [0]), .ZN(n_23_23_5));
   AOI22_X1 i_23_23_7 (.A1(\buffer[14][0][3] [0]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][3] [0]), .ZN(n_23_23_6));
   AOI22_X1 i_23_23_8 (.A1(\buffer[11][0][3] [0]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][3] [0]), .ZN(n_23_23_7));
   AOI22_X1 i_23_23_9 (.A1(\buffer[13][0][3] [0]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][3] [0]), .ZN(n_23_23_8));
   NAND4_X1 i_23_23_10 (.A1(n_23_23_17), .A2(n_23_23_15), .A3(n_23_23_13), 
      .A4(n_23_23_9), .ZN(\output_filter[0][3] [1]));
   AOI221_X1 i_23_23_11 (.A(n_23_23_10), .B1(n_25), .B2(\buffer[0][0][3] [1]), 
      .C1(\buffer[12][0][3] [1]), .C2(n_27), .ZN(n_23_23_9));
   NAND4_X1 i_23_23_12 (.A1(n_23_23_16), .A2(n_23_23_14), .A3(n_23_23_12), 
      .A4(n_23_23_11), .ZN(n_23_23_10));
   AOI22_X1 i_23_23_13 (.A1(\buffer[15][0][3] [1]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][3] [1]), .ZN(n_23_23_11));
   AOI22_X1 i_23_23_14 (.A1(\buffer[10][0][3] [1]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][3] [1]), .ZN(n_23_23_12));
   AOI22_X1 i_23_23_15 (.A1(\buffer[6][0][3] [1]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][3] [1]), .ZN(n_23_23_13));
   AOI22_X1 i_23_23_16 (.A1(\buffer[9][0][3] [1]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][3] [1]), .ZN(n_23_23_14));
   AOI22_X1 i_23_23_17 (.A1(\buffer[14][0][3] [1]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][3] [1]), .ZN(n_23_23_15));
   AOI22_X1 i_23_23_18 (.A1(\buffer[11][0][3] [1]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][3] [1]), .ZN(n_23_23_16));
   AOI22_X1 i_23_23_19 (.A1(\buffer[13][0][3] [1]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][3] [1]), .ZN(n_23_23_17));
   NAND4_X1 i_23_23_20 (.A1(n_23_23_26), .A2(n_23_23_24), .A3(n_23_23_22), 
      .A4(n_23_23_18), .ZN(\output_filter[0][3] [2]));
   AOI221_X1 i_23_23_21 (.A(n_23_23_19), .B1(n_25), .B2(\buffer[0][0][3] [2]), 
      .C1(\buffer[12][0][3] [2]), .C2(n_27), .ZN(n_23_23_18));
   NAND4_X1 i_23_23_22 (.A1(n_23_23_25), .A2(n_23_23_23), .A3(n_23_23_21), 
      .A4(n_23_23_20), .ZN(n_23_23_19));
   AOI22_X1 i_23_23_23 (.A1(\buffer[15][0][3] [2]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][3] [2]), .ZN(n_23_23_20));
   AOI22_X1 i_23_23_24 (.A1(\buffer[10][0][3] [2]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][3] [2]), .ZN(n_23_23_21));
   AOI22_X1 i_23_23_25 (.A1(\buffer[6][0][3] [2]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][3] [2]), .ZN(n_23_23_22));
   AOI22_X1 i_23_23_26 (.A1(\buffer[9][0][3] [2]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][3] [2]), .ZN(n_23_23_23));
   AOI22_X1 i_23_23_27 (.A1(\buffer[14][0][3] [2]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][3] [2]), .ZN(n_23_23_24));
   AOI22_X1 i_23_23_28 (.A1(\buffer[11][0][3] [2]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][3] [2]), .ZN(n_23_23_25));
   AOI22_X1 i_23_23_29 (.A1(\buffer[13][0][3] [2]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][3] [2]), .ZN(n_23_23_26));
   NAND4_X1 i_23_23_30 (.A1(n_23_23_35), .A2(n_23_23_33), .A3(n_23_23_31), 
      .A4(n_23_23_27), .ZN(\output_filter[0][3] [3]));
   AOI221_X1 i_23_23_31 (.A(n_23_23_28), .B1(n_25), .B2(\buffer[0][0][3] [3]), 
      .C1(\buffer[12][0][3] [3]), .C2(n_27), .ZN(n_23_23_27));
   NAND4_X1 i_23_23_32 (.A1(n_23_23_34), .A2(n_23_23_32), .A3(n_23_23_30), 
      .A4(n_23_23_29), .ZN(n_23_23_28));
   AOI22_X1 i_23_23_33 (.A1(\buffer[15][0][3] [3]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][3] [3]), .ZN(n_23_23_29));
   AOI22_X1 i_23_23_34 (.A1(\buffer[10][0][3] [3]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][3] [3]), .ZN(n_23_23_30));
   AOI22_X1 i_23_23_35 (.A1(\buffer[6][0][3] [3]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][3] [3]), .ZN(n_23_23_31));
   AOI22_X1 i_23_23_36 (.A1(\buffer[9][0][3] [3]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][3] [3]), .ZN(n_23_23_32));
   AOI22_X1 i_23_23_37 (.A1(\buffer[14][0][3] [3]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][3] [3]), .ZN(n_23_23_33));
   AOI22_X1 i_23_23_38 (.A1(\buffer[11][0][3] [3]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][3] [3]), .ZN(n_23_23_34));
   AOI22_X1 i_23_23_39 (.A1(\buffer[13][0][3] [3]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][3] [3]), .ZN(n_23_23_35));
   NAND4_X1 i_23_23_40 (.A1(n_23_23_44), .A2(n_23_23_42), .A3(n_23_23_40), 
      .A4(n_23_23_36), .ZN(\output_filter[0][3] [4]));
   AOI221_X1 i_23_23_41 (.A(n_23_23_37), .B1(n_25), .B2(\buffer[0][0][3] [4]), 
      .C1(\buffer[12][0][3] [4]), .C2(n_27), .ZN(n_23_23_36));
   NAND4_X1 i_23_23_42 (.A1(n_23_23_43), .A2(n_23_23_41), .A3(n_23_23_39), 
      .A4(n_23_23_38), .ZN(n_23_23_37));
   AOI22_X1 i_23_23_43 (.A1(\buffer[15][0][3] [4]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][3] [4]), .ZN(n_23_23_38));
   AOI22_X1 i_23_23_44 (.A1(\buffer[10][0][3] [4]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][3] [4]), .ZN(n_23_23_39));
   AOI22_X1 i_23_23_45 (.A1(\buffer[6][0][3] [4]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][3] [4]), .ZN(n_23_23_40));
   AOI22_X1 i_23_23_46 (.A1(\buffer[9][0][3] [4]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][0][3] [4]), .ZN(n_23_23_41));
   AOI22_X1 i_23_23_47 (.A1(\buffer[14][0][3] [4]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][3] [4]), .ZN(n_23_23_42));
   AOI22_X1 i_23_23_48 (.A1(\buffer[11][0][3] [4]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][3] [4]), .ZN(n_23_23_43));
   AOI22_X1 i_23_23_49 (.A1(\buffer[13][0][3] [4]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][0][3] [4]), .ZN(n_23_23_44));
   NAND4_X1 i_23_23_50 (.A1(n_23_23_53), .A2(n_23_23_51), .A3(n_23_23_49), 
      .A4(n_23_23_45), .ZN(\output_filter[0][3] [5]));
   AOI221_X1 i_23_23_51 (.A(n_23_23_46), .B1(n_25), .B2(\buffer[0][0][3] [5]), 
      .C1(\buffer[12][0][3] [5]), .C2(n_27), .ZN(n_23_23_45));
   NAND4_X1 i_23_23_52 (.A1(n_23_23_52), .A2(n_23_23_50), .A3(n_23_23_48), 
      .A4(n_23_23_47), .ZN(n_23_23_46));
   AOI22_X1 i_23_23_53 (.A1(\buffer[15][0][3] [5]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][3] [5]), .ZN(n_23_23_47));
   AOI22_X1 i_23_23_54 (.A1(\buffer[10][0][3] [5]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][3] [5]), .ZN(n_23_23_48));
   AOI22_X1 i_23_23_55 (.A1(\buffer[6][0][3] [5]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][3] [5]), .ZN(n_23_23_49));
   AOI22_X1 i_23_23_56 (.A1(\buffer[9][0][3] [5]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][3] [5]), .ZN(n_23_23_50));
   AOI22_X1 i_23_23_57 (.A1(\buffer[14][0][3] [5]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][3] [5]), .ZN(n_23_23_51));
   AOI22_X1 i_23_23_58 (.A1(\buffer[11][0][3] [5]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][3] [5]), .ZN(n_23_23_52));
   AOI22_X1 i_23_23_59 (.A1(\buffer[13][0][3] [5]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][3] [5]), .ZN(n_23_23_53));
   NAND4_X1 i_23_23_60 (.A1(n_23_23_62), .A2(n_23_23_60), .A3(n_23_23_58), 
      .A4(n_23_23_54), .ZN(\output_filter[0][3] [6]));
   AOI221_X1 i_23_23_61 (.A(n_23_23_55), .B1(n_25), .B2(\buffer[0][0][3] [6]), 
      .C1(\buffer[12][0][3] [6]), .C2(n_27), .ZN(n_23_23_54));
   NAND4_X1 i_23_23_62 (.A1(n_23_23_61), .A2(n_23_23_59), .A3(n_23_23_57), 
      .A4(n_23_23_56), .ZN(n_23_23_55));
   AOI22_X1 i_23_23_63 (.A1(\buffer[15][0][3] [6]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][3] [6]), .ZN(n_23_23_56));
   AOI22_X1 i_23_23_64 (.A1(\buffer[10][0][3] [6]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][3] [6]), .ZN(n_23_23_57));
   AOI22_X1 i_23_23_65 (.A1(\buffer[6][0][3] [6]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][3] [6]), .ZN(n_23_23_58));
   AOI22_X1 i_23_23_66 (.A1(\buffer[9][0][3] [6]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][3] [6]), .ZN(n_23_23_59));
   AOI22_X1 i_23_23_67 (.A1(\buffer[14][0][3] [6]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][3] [6]), .ZN(n_23_23_60));
   AOI22_X1 i_23_23_68 (.A1(\buffer[11][0][3] [6]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][3] [6]), .ZN(n_23_23_61));
   AOI22_X1 i_23_23_69 (.A1(\buffer[13][0][3] [6]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][3] [6]), .ZN(n_23_23_62));
   NAND4_X1 i_23_23_70 (.A1(n_23_23_71), .A2(n_23_23_69), .A3(n_23_23_67), 
      .A4(n_23_23_63), .ZN(\output_filter[0][3] [7]));
   AOI221_X1 i_23_23_71 (.A(n_23_23_64), .B1(n_25), .B2(\buffer[0][0][3] [7]), 
      .C1(\buffer[12][0][3] [7]), .C2(n_27), .ZN(n_23_23_63));
   NAND4_X1 i_23_23_72 (.A1(n_23_23_70), .A2(n_23_23_68), .A3(n_23_23_66), 
      .A4(n_23_23_65), .ZN(n_23_23_64));
   AOI22_X1 i_23_23_73 (.A1(\buffer[15][0][3] [7]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][3] [7]), .ZN(n_23_23_65));
   AOI22_X1 i_23_23_74 (.A1(\buffer[10][0][3] [7]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][3] [7]), .ZN(n_23_23_66));
   AOI22_X1 i_23_23_75 (.A1(\buffer[6][0][3] [7]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][3] [7]), .ZN(n_23_23_67));
   AOI22_X1 i_23_23_76 (.A1(\buffer[9][0][3] [7]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][0][3] [7]), .ZN(n_23_23_68));
   AOI22_X1 i_23_23_77 (.A1(\buffer[14][0][3] [7]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][3] [7]), .ZN(n_23_23_69));
   AOI22_X1 i_23_23_78 (.A1(\buffer[11][0][3] [7]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][3] [7]), .ZN(n_23_23_70));
   AOI22_X1 i_23_23_79 (.A1(\buffer[13][0][3] [7]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][0][3] [7]), .ZN(n_23_23_71));
   NAND4_X1 i_23_23_80 (.A1(n_23_23_80), .A2(n_23_23_78), .A3(n_23_23_76), 
      .A4(n_23_23_72), .ZN(\output_filter[0][3] [8]));
   AOI221_X1 i_23_23_81 (.A(n_23_23_73), .B1(n_25), .B2(\buffer[0][0][3] [8]), 
      .C1(\buffer[12][0][3] [8]), .C2(n_27), .ZN(n_23_23_72));
   NAND4_X1 i_23_23_82 (.A1(n_23_23_79), .A2(n_23_23_77), .A3(n_23_23_75), 
      .A4(n_23_23_74), .ZN(n_23_23_73));
   AOI22_X1 i_23_23_83 (.A1(\buffer[15][0][3] [8]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][3] [8]), .ZN(n_23_23_74));
   AOI22_X1 i_23_23_84 (.A1(\buffer[10][0][3] [8]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][3] [8]), .ZN(n_23_23_75));
   AOI22_X1 i_23_23_85 (.A1(\buffer[6][0][3] [8]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][3] [8]), .ZN(n_23_23_76));
   AOI22_X1 i_23_23_86 (.A1(\buffer[9][0][3] [8]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][3] [8]), .ZN(n_23_23_77));
   AOI22_X1 i_23_23_87 (.A1(\buffer[14][0][3] [8]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][3] [8]), .ZN(n_23_23_78));
   AOI22_X1 i_23_23_88 (.A1(\buffer[11][0][3] [8]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][3] [8]), .ZN(n_23_23_79));
   AOI22_X1 i_23_23_89 (.A1(\buffer[13][0][3] [8]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][3] [8]), .ZN(n_23_23_80));
   NAND4_X1 i_23_23_90 (.A1(n_23_23_89), .A2(n_23_23_87), .A3(n_23_23_85), 
      .A4(n_23_23_81), .ZN(\output_filter[0][3] [9]));
   AOI221_X1 i_23_23_91 (.A(n_23_23_82), .B1(n_25), .B2(\buffer[0][0][3] [9]), 
      .C1(\buffer[12][0][3] [9]), .C2(n_27), .ZN(n_23_23_81));
   NAND4_X1 i_23_23_92 (.A1(n_23_23_88), .A2(n_23_23_86), .A3(n_23_23_84), 
      .A4(n_23_23_83), .ZN(n_23_23_82));
   AOI22_X1 i_23_23_93 (.A1(\buffer[15][0][3] [9]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][3] [9]), .ZN(n_23_23_83));
   AOI22_X1 i_23_23_94 (.A1(\buffer[10][0][3] [9]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][3] [9]), .ZN(n_23_23_84));
   AOI22_X1 i_23_23_95 (.A1(\buffer[6][0][3] [9]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][3] [9]), .ZN(n_23_23_85));
   AOI22_X1 i_23_23_96 (.A1(\buffer[9][0][3] [9]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][0][3] [9]), .ZN(n_23_23_86));
   AOI22_X1 i_23_23_97 (.A1(\buffer[14][0][3] [9]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][3] [9]), .ZN(n_23_23_87));
   AOI22_X1 i_23_23_98 (.A1(\buffer[11][0][3] [9]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][3] [9]), .ZN(n_23_23_88));
   AOI22_X1 i_23_23_99 (.A1(\buffer[13][0][3] [9]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][0][3] [9]), .ZN(n_23_23_89));
   NAND4_X1 i_23_23_100 (.A1(n_23_23_98), .A2(n_23_23_96), .A3(n_23_23_94), 
      .A4(n_23_23_90), .ZN(\output_filter[0][3] [10]));
   AOI221_X1 i_23_23_101 (.A(n_23_23_91), .B1(n_25), .B2(\buffer[0][0][3] [10]), 
      .C1(\buffer[12][0][3] [10]), .C2(n_27), .ZN(n_23_23_90));
   NAND4_X1 i_23_23_102 (.A1(n_23_23_97), .A2(n_23_23_95), .A3(n_23_23_93), 
      .A4(n_23_23_92), .ZN(n_23_23_91));
   AOI22_X1 i_23_23_103 (.A1(\buffer[15][0][3] [10]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][3] [10]), .ZN(n_23_23_92));
   AOI22_X1 i_23_23_104 (.A1(\buffer[10][0][3] [10]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][3] [10]), .ZN(n_23_23_93));
   AOI22_X1 i_23_23_105 (.A1(\buffer[6][0][3] [10]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][3] [10]), .ZN(n_23_23_94));
   AOI22_X1 i_23_23_106 (.A1(\buffer[9][0][3] [10]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][3] [10]), .ZN(n_23_23_95));
   AOI22_X1 i_23_23_107 (.A1(\buffer[14][0][3] [10]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][3] [10]), .ZN(n_23_23_96));
   AOI22_X1 i_23_23_108 (.A1(\buffer[11][0][3] [10]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][3] [10]), .ZN(n_23_23_97));
   AOI22_X1 i_23_23_109 (.A1(\buffer[13][0][3] [10]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][3] [10]), .ZN(n_23_23_98));
   NAND4_X1 i_23_23_110 (.A1(n_23_23_107), .A2(n_23_23_105), .A3(n_23_23_103), 
      .A4(n_23_23_99), .ZN(\output_filter[0][3] [11]));
   AOI221_X1 i_23_23_111 (.A(n_23_23_100), .B1(n_25), .B2(\buffer[0][0][3] [11]), 
      .C1(\buffer[12][0][3] [11]), .C2(n_27), .ZN(n_23_23_99));
   NAND4_X1 i_23_23_112 (.A1(n_23_23_106), .A2(n_23_23_104), .A3(n_23_23_102), 
      .A4(n_23_23_101), .ZN(n_23_23_100));
   AOI22_X1 i_23_23_113 (.A1(\buffer[15][0][3] [11]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][3] [11]), .ZN(n_23_23_101));
   AOI22_X1 i_23_23_114 (.A1(\buffer[10][0][3] [11]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][3] [11]), .ZN(n_23_23_102));
   AOI22_X1 i_23_23_115 (.A1(\buffer[6][0][3] [11]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][3] [11]), .ZN(n_23_23_103));
   AOI22_X1 i_23_23_116 (.A1(\buffer[9][0][3] [11]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][0][3] [11]), .ZN(n_23_23_104));
   AOI22_X1 i_23_23_117 (.A1(\buffer[14][0][3] [11]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][3] [11]), .ZN(n_23_23_105));
   AOI22_X1 i_23_23_118 (.A1(\buffer[11][0][3] [11]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][3] [11]), .ZN(n_23_23_106));
   AOI22_X1 i_23_23_119 (.A1(\buffer[13][0][3] [11]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][0][3] [11]), .ZN(n_23_23_107));
   NAND4_X1 i_23_23_120 (.A1(n_23_23_116), .A2(n_23_23_114), .A3(n_23_23_112), 
      .A4(n_23_23_108), .ZN(\output_filter[0][3] [12]));
   AOI221_X1 i_23_23_121 (.A(n_23_23_109), .B1(n_25), .B2(\buffer[0][0][3] [12]), 
      .C1(\buffer[12][0][3] [12]), .C2(n_27), .ZN(n_23_23_108));
   NAND4_X1 i_23_23_122 (.A1(n_23_23_115), .A2(n_23_23_113), .A3(n_23_23_111), 
      .A4(n_23_23_110), .ZN(n_23_23_109));
   AOI22_X1 i_23_23_123 (.A1(\buffer[15][0][3] [12]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][3] [12]), .ZN(n_23_23_110));
   AOI22_X1 i_23_23_124 (.A1(\buffer[10][0][3] [12]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][3] [12]), .ZN(n_23_23_111));
   AOI22_X1 i_23_23_125 (.A1(\buffer[6][0][3] [12]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][3] [12]), .ZN(n_23_23_112));
   AOI22_X1 i_23_23_126 (.A1(\buffer[9][0][3] [12]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][3] [12]), .ZN(n_23_23_113));
   AOI22_X1 i_23_23_127 (.A1(\buffer[14][0][3] [12]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][3] [12]), .ZN(n_23_23_114));
   AOI22_X1 i_23_23_128 (.A1(\buffer[11][0][3] [12]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][3] [12]), .ZN(n_23_23_115));
   AOI22_X1 i_23_23_129 (.A1(\buffer[13][0][3] [12]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][3] [12]), .ZN(n_23_23_116));
   NAND4_X1 i_23_23_130 (.A1(n_23_23_125), .A2(n_23_23_123), .A3(n_23_23_121), 
      .A4(n_23_23_117), .ZN(\output_filter[0][3] [13]));
   AOI221_X1 i_23_23_131 (.A(n_23_23_118), .B1(n_25), .B2(\buffer[0][0][3] [13]), 
      .C1(\buffer[12][0][3] [13]), .C2(n_27), .ZN(n_23_23_117));
   NAND4_X1 i_23_23_132 (.A1(n_23_23_124), .A2(n_23_23_122), .A3(n_23_23_120), 
      .A4(n_23_23_119), .ZN(n_23_23_118));
   AOI22_X1 i_23_23_133 (.A1(\buffer[15][0][3] [13]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][3] [13]), .ZN(n_23_23_119));
   AOI22_X1 i_23_23_134 (.A1(\buffer[10][0][3] [13]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][3] [13]), .ZN(n_23_23_120));
   AOI22_X1 i_23_23_135 (.A1(\buffer[6][0][3] [13]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][3] [13]), .ZN(n_23_23_121));
   AOI22_X1 i_23_23_136 (.A1(\buffer[9][0][3] [13]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][0][3] [13]), .ZN(n_23_23_122));
   AOI22_X1 i_23_23_137 (.A1(\buffer[14][0][3] [13]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][3] [13]), .ZN(n_23_23_123));
   AOI22_X1 i_23_23_138 (.A1(\buffer[11][0][3] [13]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][3] [13]), .ZN(n_23_23_124));
   AOI22_X1 i_23_23_139 (.A1(\buffer[13][0][3] [13]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][0][3] [13]), .ZN(n_23_23_125));
   NAND4_X1 i_23_23_140 (.A1(n_23_23_134), .A2(n_23_23_132), .A3(n_23_23_130), 
      .A4(n_23_23_126), .ZN(\output_filter[0][3] [14]));
   AOI221_X1 i_23_23_141 (.A(n_23_23_127), .B1(n_25), .B2(\buffer[0][0][3] [14]), 
      .C1(\buffer[12][0][3] [14]), .C2(n_27), .ZN(n_23_23_126));
   NAND4_X1 i_23_23_142 (.A1(n_23_23_133), .A2(n_23_23_131), .A3(n_23_23_129), 
      .A4(n_23_23_128), .ZN(n_23_23_127));
   AOI22_X1 i_23_23_143 (.A1(\buffer[15][0][3] [14]), .A2(n_22), .B1(n_16), 
      .B2(\buffer[8][0][3] [14]), .ZN(n_23_23_128));
   AOI22_X1 i_23_23_144 (.A1(\buffer[10][0][3] [14]), .A2(n_21), .B1(n_29), 
      .B2(\buffer[7][0][3] [14]), .ZN(n_23_23_129));
   AOI22_X1 i_23_23_145 (.A1(\buffer[6][0][3] [14]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][3] [14]), .ZN(n_23_23_130));
   AOI22_X1 i_23_23_146 (.A1(\buffer[9][0][3] [14]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][3] [14]), .ZN(n_23_23_131));
   AOI22_X1 i_23_23_147 (.A1(\buffer[14][0][3] [14]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][3] [14]), .ZN(n_23_23_132));
   AOI22_X1 i_23_23_148 (.A1(\buffer[11][0][3] [14]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][3] [14]), .ZN(n_23_23_133));
   AOI22_X1 i_23_23_149 (.A1(\buffer[13][0][3] [14]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][3] [14]), .ZN(n_23_23_134));
   NAND2_X1 i_23_23_150 (.A1(n_23_23_137), .A2(n_23_23_135), .ZN(
      \output_filter[0][3] [15]));
   AOI221_X1 i_23_23_151 (.A(n_23_23_136), .B1(n_31), .B2(\buffer[3][0][3] [15]), 
      .C1(\buffer[14][0][3] [15]), .C2(n_19), .ZN(n_23_23_135));
   NAND3_X1 i_23_23_152 (.A1(n_23_23_143), .A2(n_23_23_141), .A3(n_23_23_139), 
      .ZN(n_23_23_136));
   AOI221_X1 i_23_23_153 (.A(n_23_23_138), .B1(n_16), .B2(\buffer[8][0][3] [15]), 
      .C1(\buffer[13][0][3] [15]), .C2(n_26), .ZN(n_23_23_137));
   NAND3_X1 i_23_23_154 (.A1(n_23_23_144), .A2(n_23_23_142), .A3(n_23_23_140), 
      .ZN(n_23_23_138));
   AOI22_X1 i_23_23_155 (.A1(\buffer[11][0][3] [15]), .A2(n_17), .B1(n_24), 
      .B2(\buffer[2][0][3] [15]), .ZN(n_23_23_139));
   AOI22_X1 i_23_23_156 (.A1(\buffer[10][0][3] [15]), .A2(n_21), .B1(n_23), 
      .B2(\buffer[1][0][3] [15]), .ZN(n_23_23_140));
   AOI22_X1 i_23_23_157 (.A1(\buffer[6][0][3] [15]), .A2(n_28), .B1(n_18), 
      .B2(\buffer[5][0][3] [15]), .ZN(n_23_23_141));
   AOI22_X1 i_23_23_158 (.A1(\buffer[9][0][3] [15]), .A2(n_20), .B1(n_30), 
      .B2(\buffer[4][0][3] [15]), .ZN(n_23_23_142));
   AOI22_X1 i_23_23_159 (.A1(\buffer[7][0][3] [15]), .A2(n_29), .B1(n_25), 
      .B2(\buffer[0][0][3] [15]), .ZN(n_23_23_143));
   AOI22_X1 i_23_23_160 (.A1(\buffer[15][0][3] [15]), .A2(n_22), .B1(n_27), 
      .B2(\buffer[12][0][3] [15]), .ZN(n_23_23_144));
   NAND4_X1 i_22_22_0 (.A1(n_22_22_8), .A2(n_22_22_6), .A3(n_22_22_4), .A4(
      n_22_22_0), .ZN(\output_filter[0][2] [0]));
   AOI221_X1 i_22_22_1 (.A(n_22_22_1), .B1(n_25), .B2(\buffer[0][0][2] [0]), 
      .C1(\buffer[12][0][2] [0]), .C2(n_27), .ZN(n_22_22_0));
   NAND4_X1 i_22_22_2 (.A1(n_22_22_7), .A2(n_22_22_5), .A3(n_22_22_3), .A4(
      n_22_22_2), .ZN(n_22_22_1));
   AOI22_X1 i_22_22_3 (.A1(\buffer[15][0][2] [0]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][2] [0]), .ZN(n_22_22_2));
   AOI22_X1 i_22_22_4 (.A1(\buffer[10][0][2] [0]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][2] [0]), .ZN(n_22_22_3));
   AOI22_X1 i_22_22_5 (.A1(\buffer[6][0][2] [0]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][0][2] [0]), .ZN(n_22_22_4));
   AOI22_X1 i_22_22_6 (.A1(\buffer[9][0][2] [0]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][0][2] [0]), .ZN(n_22_22_5));
   AOI22_X1 i_22_22_7 (.A1(\buffer[14][0][2] [0]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][2] [0]), .ZN(n_22_22_6));
   AOI22_X1 i_22_22_8 (.A1(\buffer[11][0][2] [0]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][2] [0]), .ZN(n_22_22_7));
   AOI22_X1 i_22_22_9 (.A1(\buffer[13][0][2] [0]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][2] [0]), .ZN(n_22_22_8));
   NAND4_X1 i_22_22_10 (.A1(n_22_22_17), .A2(n_22_22_15), .A3(n_22_22_13), 
      .A4(n_22_22_9), .ZN(\output_filter[0][2] [1]));
   AOI221_X1 i_22_22_11 (.A(n_22_22_10), .B1(n_25), .B2(\buffer[0][0][2] [1]), 
      .C1(\buffer[12][0][2] [1]), .C2(n_27), .ZN(n_22_22_9));
   NAND4_X1 i_22_22_12 (.A1(n_22_22_16), .A2(n_22_22_14), .A3(n_22_22_12), 
      .A4(n_22_22_11), .ZN(n_22_22_10));
   AOI22_X1 i_22_22_13 (.A1(\buffer[15][0][2] [1]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][2] [1]), .ZN(n_22_22_11));
   AOI22_X1 i_22_22_14 (.A1(\buffer[10][0][2] [1]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][2] [1]), .ZN(n_22_22_12));
   AOI22_X1 i_22_22_15 (.A1(\buffer[6][0][2] [1]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][2] [1]), .ZN(n_22_22_13));
   AOI22_X1 i_22_22_16 (.A1(\buffer[9][0][2] [1]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][2] [1]), .ZN(n_22_22_14));
   AOI22_X1 i_22_22_17 (.A1(\buffer[14][0][2] [1]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][2] [1]), .ZN(n_22_22_15));
   AOI22_X1 i_22_22_18 (.A1(\buffer[11][0][2] [1]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][2] [1]), .ZN(n_22_22_16));
   AOI22_X1 i_22_22_19 (.A1(\buffer[13][0][2] [1]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][2] [1]), .ZN(n_22_22_17));
   NAND4_X1 i_22_22_20 (.A1(n_22_22_26), .A2(n_22_22_24), .A3(n_22_22_22), 
      .A4(n_22_22_18), .ZN(\output_filter[0][2] [2]));
   AOI221_X1 i_22_22_21 (.A(n_22_22_19), .B1(n_25), .B2(\buffer[0][0][2] [2]), 
      .C1(\buffer[12][0][2] [2]), .C2(n_27), .ZN(n_22_22_18));
   NAND4_X1 i_22_22_22 (.A1(n_22_22_25), .A2(n_22_22_23), .A3(n_22_22_21), 
      .A4(n_22_22_20), .ZN(n_22_22_19));
   AOI22_X1 i_22_22_23 (.A1(\buffer[15][0][2] [2]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][2] [2]), .ZN(n_22_22_20));
   AOI22_X1 i_22_22_24 (.A1(\buffer[10][0][2] [2]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][2] [2]), .ZN(n_22_22_21));
   AOI22_X1 i_22_22_25 (.A1(\buffer[6][0][2] [2]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][2] [2]), .ZN(n_22_22_22));
   AOI22_X1 i_22_22_26 (.A1(\buffer[9][0][2] [2]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][2] [2]), .ZN(n_22_22_23));
   AOI22_X1 i_22_22_27 (.A1(\buffer[14][0][2] [2]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][2] [2]), .ZN(n_22_22_24));
   AOI22_X1 i_22_22_28 (.A1(\buffer[11][0][2] [2]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][2] [2]), .ZN(n_22_22_25));
   AOI22_X1 i_22_22_29 (.A1(\buffer[13][0][2] [2]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][2] [2]), .ZN(n_22_22_26));
   NAND4_X1 i_22_22_30 (.A1(n_22_22_35), .A2(n_22_22_33), .A3(n_22_22_31), 
      .A4(n_22_22_27), .ZN(\output_filter[0][2] [3]));
   AOI221_X1 i_22_22_31 (.A(n_22_22_28), .B1(n_25), .B2(\buffer[0][0][2] [3]), 
      .C1(\buffer[12][0][2] [3]), .C2(n_27), .ZN(n_22_22_27));
   NAND4_X1 i_22_22_32 (.A1(n_22_22_34), .A2(n_22_22_32), .A3(n_22_22_30), 
      .A4(n_22_22_29), .ZN(n_22_22_28));
   AOI22_X1 i_22_22_33 (.A1(\buffer[15][0][2] [3]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][2] [3]), .ZN(n_22_22_29));
   AOI22_X1 i_22_22_34 (.A1(\buffer[10][0][2] [3]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][2] [3]), .ZN(n_22_22_30));
   AOI22_X1 i_22_22_35 (.A1(\buffer[6][0][2] [3]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][2] [3]), .ZN(n_22_22_31));
   AOI22_X1 i_22_22_36 (.A1(\buffer[9][0][2] [3]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][2] [3]), .ZN(n_22_22_32));
   AOI22_X1 i_22_22_37 (.A1(\buffer[14][0][2] [3]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][2] [3]), .ZN(n_22_22_33));
   AOI22_X1 i_22_22_38 (.A1(\buffer[11][0][2] [3]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][2] [3]), .ZN(n_22_22_34));
   AOI22_X1 i_22_22_39 (.A1(\buffer[13][0][2] [3]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][2] [3]), .ZN(n_22_22_35));
   NAND4_X1 i_22_22_40 (.A1(n_22_22_44), .A2(n_22_22_42), .A3(n_22_22_40), 
      .A4(n_22_22_36), .ZN(\output_filter[0][2] [4]));
   AOI221_X1 i_22_22_41 (.A(n_22_22_37), .B1(n_25), .B2(\buffer[0][0][2] [4]), 
      .C1(\buffer[12][0][2] [4]), .C2(n_27), .ZN(n_22_22_36));
   NAND4_X1 i_22_22_42 (.A1(n_22_22_43), .A2(n_22_22_41), .A3(n_22_22_39), 
      .A4(n_22_22_38), .ZN(n_22_22_37));
   AOI22_X1 i_22_22_43 (.A1(\buffer[15][0][2] [4]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][2] [4]), .ZN(n_22_22_38));
   AOI22_X1 i_22_22_44 (.A1(\buffer[10][0][2] [4]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][2] [4]), .ZN(n_22_22_39));
   AOI22_X1 i_22_22_45 (.A1(\buffer[6][0][2] [4]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][2] [4]), .ZN(n_22_22_40));
   AOI22_X1 i_22_22_46 (.A1(\buffer[9][0][2] [4]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][0][2] [4]), .ZN(n_22_22_41));
   AOI22_X1 i_22_22_47 (.A1(\buffer[14][0][2] [4]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][2] [4]), .ZN(n_22_22_42));
   AOI22_X1 i_22_22_48 (.A1(\buffer[11][0][2] [4]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][2] [4]), .ZN(n_22_22_43));
   AOI22_X1 i_22_22_49 (.A1(\buffer[13][0][2] [4]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][0][2] [4]), .ZN(n_22_22_44));
   NAND4_X1 i_22_22_50 (.A1(n_22_22_53), .A2(n_22_22_51), .A3(n_22_22_49), 
      .A4(n_22_22_45), .ZN(\output_filter[0][2] [5]));
   AOI221_X1 i_22_22_51 (.A(n_22_22_46), .B1(n_25), .B2(\buffer[0][0][2] [5]), 
      .C1(\buffer[12][0][2] [5]), .C2(n_27), .ZN(n_22_22_45));
   NAND4_X1 i_22_22_52 (.A1(n_22_22_52), .A2(n_22_22_50), .A3(n_22_22_48), 
      .A4(n_22_22_47), .ZN(n_22_22_46));
   AOI22_X1 i_22_22_53 (.A1(\buffer[15][0][2] [5]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][2] [5]), .ZN(n_22_22_47));
   AOI22_X1 i_22_22_54 (.A1(\buffer[10][0][2] [5]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][2] [5]), .ZN(n_22_22_48));
   AOI22_X1 i_22_22_55 (.A1(\buffer[6][0][2] [5]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][2] [5]), .ZN(n_22_22_49));
   AOI22_X1 i_22_22_56 (.A1(\buffer[9][0][2] [5]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][2] [5]), .ZN(n_22_22_50));
   AOI22_X1 i_22_22_57 (.A1(\buffer[14][0][2] [5]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][2] [5]), .ZN(n_22_22_51));
   AOI22_X1 i_22_22_58 (.A1(\buffer[11][0][2] [5]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][2] [5]), .ZN(n_22_22_52));
   AOI22_X1 i_22_22_59 (.A1(\buffer[13][0][2] [5]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][2] [5]), .ZN(n_22_22_53));
   NAND4_X1 i_22_22_60 (.A1(n_22_22_62), .A2(n_22_22_60), .A3(n_22_22_58), 
      .A4(n_22_22_54), .ZN(\output_filter[0][2] [6]));
   AOI221_X1 i_22_22_61 (.A(n_22_22_55), .B1(n_25), .B2(\buffer[0][0][2] [6]), 
      .C1(\buffer[12][0][2] [6]), .C2(n_27), .ZN(n_22_22_54));
   NAND4_X1 i_22_22_62 (.A1(n_22_22_61), .A2(n_22_22_59), .A3(n_22_22_57), 
      .A4(n_22_22_56), .ZN(n_22_22_55));
   AOI22_X1 i_22_22_63 (.A1(\buffer[15][0][2] [6]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][2] [6]), .ZN(n_22_22_56));
   AOI22_X1 i_22_22_64 (.A1(\buffer[10][0][2] [6]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][2] [6]), .ZN(n_22_22_57));
   AOI22_X1 i_22_22_65 (.A1(\buffer[6][0][2] [6]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][2] [6]), .ZN(n_22_22_58));
   AOI22_X1 i_22_22_66 (.A1(\buffer[9][0][2] [6]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][2] [6]), .ZN(n_22_22_59));
   AOI22_X1 i_22_22_67 (.A1(\buffer[14][0][2] [6]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][2] [6]), .ZN(n_22_22_60));
   AOI22_X1 i_22_22_68 (.A1(\buffer[11][0][2] [6]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][2] [6]), .ZN(n_22_22_61));
   AOI22_X1 i_22_22_69 (.A1(\buffer[13][0][2] [6]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][2] [6]), .ZN(n_22_22_62));
   NAND4_X1 i_22_22_70 (.A1(n_22_22_71), .A2(n_22_22_69), .A3(n_22_22_67), 
      .A4(n_22_22_63), .ZN(\output_filter[0][2] [7]));
   AOI221_X1 i_22_22_71 (.A(n_22_22_64), .B1(n_25), .B2(\buffer[0][0][2] [7]), 
      .C1(\buffer[12][0][2] [7]), .C2(n_27), .ZN(n_22_22_63));
   NAND4_X1 i_22_22_72 (.A1(n_22_22_70), .A2(n_22_22_68), .A3(n_22_22_66), 
      .A4(n_22_22_65), .ZN(n_22_22_64));
   AOI22_X1 i_22_22_73 (.A1(\buffer[15][0][2] [7]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][2] [7]), .ZN(n_22_22_65));
   AOI22_X1 i_22_22_74 (.A1(\buffer[10][0][2] [7]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][2] [7]), .ZN(n_22_22_66));
   AOI22_X1 i_22_22_75 (.A1(\buffer[6][0][2] [7]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][2] [7]), .ZN(n_22_22_67));
   AOI22_X1 i_22_22_76 (.A1(\buffer[9][0][2] [7]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][0][2] [7]), .ZN(n_22_22_68));
   AOI22_X1 i_22_22_77 (.A1(\buffer[14][0][2] [7]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][2] [7]), .ZN(n_22_22_69));
   AOI22_X1 i_22_22_78 (.A1(\buffer[11][0][2] [7]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][2] [7]), .ZN(n_22_22_70));
   AOI22_X1 i_22_22_79 (.A1(\buffer[13][0][2] [7]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][0][2] [7]), .ZN(n_22_22_71));
   NAND4_X1 i_22_22_80 (.A1(n_22_22_80), .A2(n_22_22_78), .A3(n_22_22_76), 
      .A4(n_22_22_72), .ZN(\output_filter[0][2] [8]));
   AOI221_X1 i_22_22_81 (.A(n_22_22_73), .B1(n_25), .B2(\buffer[0][0][2] [8]), 
      .C1(\buffer[12][0][2] [8]), .C2(n_27), .ZN(n_22_22_72));
   NAND4_X1 i_22_22_82 (.A1(n_22_22_79), .A2(n_22_22_77), .A3(n_22_22_75), 
      .A4(n_22_22_74), .ZN(n_22_22_73));
   AOI22_X1 i_22_22_83 (.A1(\buffer[15][0][2] [8]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][2] [8]), .ZN(n_22_22_74));
   AOI22_X1 i_22_22_84 (.A1(\buffer[10][0][2] [8]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][2] [8]), .ZN(n_22_22_75));
   AOI22_X1 i_22_22_85 (.A1(\buffer[6][0][2] [8]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][2] [8]), .ZN(n_22_22_76));
   AOI22_X1 i_22_22_86 (.A1(\buffer[9][0][2] [8]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][2] [8]), .ZN(n_22_22_77));
   AOI22_X1 i_22_22_87 (.A1(\buffer[14][0][2] [8]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][2] [8]), .ZN(n_22_22_78));
   AOI22_X1 i_22_22_88 (.A1(\buffer[11][0][2] [8]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][2] [8]), .ZN(n_22_22_79));
   AOI22_X1 i_22_22_89 (.A1(\buffer[13][0][2] [8]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][2] [8]), .ZN(n_22_22_80));
   NAND4_X1 i_22_22_90 (.A1(n_22_22_89), .A2(n_22_22_87), .A3(n_22_22_85), 
      .A4(n_22_22_81), .ZN(\output_filter[0][2] [9]));
   AOI221_X1 i_22_22_91 (.A(n_22_22_82), .B1(n_25), .B2(\buffer[0][0][2] [9]), 
      .C1(\buffer[12][0][2] [9]), .C2(n_27), .ZN(n_22_22_81));
   NAND4_X1 i_22_22_92 (.A1(n_22_22_88), .A2(n_22_22_86), .A3(n_22_22_84), 
      .A4(n_22_22_83), .ZN(n_22_22_82));
   AOI22_X1 i_22_22_93 (.A1(\buffer[15][0][2] [9]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][2] [9]), .ZN(n_22_22_83));
   AOI22_X1 i_22_22_94 (.A1(\buffer[10][0][2] [9]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][2] [9]), .ZN(n_22_22_84));
   AOI22_X1 i_22_22_95 (.A1(\buffer[6][0][2] [9]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][2] [9]), .ZN(n_22_22_85));
   AOI22_X1 i_22_22_96 (.A1(\buffer[9][0][2] [9]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][0][2] [9]), .ZN(n_22_22_86));
   AOI22_X1 i_22_22_97 (.A1(\buffer[14][0][2] [9]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][2] [9]), .ZN(n_22_22_87));
   AOI22_X1 i_22_22_98 (.A1(\buffer[11][0][2] [9]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][2] [9]), .ZN(n_22_22_88));
   AOI22_X1 i_22_22_99 (.A1(\buffer[13][0][2] [9]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][0][2] [9]), .ZN(n_22_22_89));
   NAND4_X1 i_22_22_100 (.A1(n_22_22_98), .A2(n_22_22_96), .A3(n_22_22_94), 
      .A4(n_22_22_90), .ZN(\output_filter[0][2] [10]));
   AOI221_X1 i_22_22_101 (.A(n_22_22_91), .B1(n_25), .B2(\buffer[0][0][2] [10]), 
      .C1(\buffer[12][0][2] [10]), .C2(n_27), .ZN(n_22_22_90));
   NAND4_X1 i_22_22_102 (.A1(n_22_22_97), .A2(n_22_22_95), .A3(n_22_22_93), 
      .A4(n_22_22_92), .ZN(n_22_22_91));
   AOI22_X1 i_22_22_103 (.A1(\buffer[15][0][2] [10]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][2] [10]), .ZN(n_22_22_92));
   AOI22_X1 i_22_22_104 (.A1(\buffer[10][0][2] [10]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][2] [10]), .ZN(n_22_22_93));
   AOI22_X1 i_22_22_105 (.A1(\buffer[6][0][2] [10]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][2] [10]), .ZN(n_22_22_94));
   AOI22_X1 i_22_22_106 (.A1(\buffer[9][0][2] [10]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][2] [10]), .ZN(n_22_22_95));
   AOI22_X1 i_22_22_107 (.A1(\buffer[14][0][2] [10]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][2] [10]), .ZN(n_22_22_96));
   AOI22_X1 i_22_22_108 (.A1(\buffer[11][0][2] [10]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][2] [10]), .ZN(n_22_22_97));
   AOI22_X1 i_22_22_109 (.A1(\buffer[13][0][2] [10]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][2] [10]), .ZN(n_22_22_98));
   NAND4_X1 i_22_22_110 (.A1(n_22_22_107), .A2(n_22_22_105), .A3(n_22_22_103), 
      .A4(n_22_22_99), .ZN(\output_filter[0][2] [11]));
   AOI221_X1 i_22_22_111 (.A(n_22_22_100), .B1(n_25), .B2(\buffer[0][0][2] [11]), 
      .C1(\buffer[12][0][2] [11]), .C2(n_27), .ZN(n_22_22_99));
   NAND4_X1 i_22_22_112 (.A1(n_22_22_106), .A2(n_22_22_104), .A3(n_22_22_102), 
      .A4(n_22_22_101), .ZN(n_22_22_100));
   AOI22_X1 i_22_22_113 (.A1(\buffer[15][0][2] [11]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][2] [11]), .ZN(n_22_22_101));
   AOI22_X1 i_22_22_114 (.A1(\buffer[10][0][2] [11]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][2] [11]), .ZN(n_22_22_102));
   AOI22_X1 i_22_22_115 (.A1(\buffer[6][0][2] [11]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][2] [11]), .ZN(n_22_22_103));
   AOI22_X1 i_22_22_116 (.A1(\buffer[9][0][2] [11]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][0][2] [11]), .ZN(n_22_22_104));
   AOI22_X1 i_22_22_117 (.A1(\buffer[14][0][2] [11]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][2] [11]), .ZN(n_22_22_105));
   AOI22_X1 i_22_22_118 (.A1(\buffer[11][0][2] [11]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][2] [11]), .ZN(n_22_22_106));
   AOI22_X1 i_22_22_119 (.A1(\buffer[13][0][2] [11]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][0][2] [11]), .ZN(n_22_22_107));
   NAND4_X1 i_22_22_120 (.A1(n_22_22_116), .A2(n_22_22_114), .A3(n_22_22_112), 
      .A4(n_22_22_108), .ZN(\output_filter[0][2] [12]));
   AOI221_X1 i_22_22_121 (.A(n_22_22_109), .B1(n_25), .B2(\buffer[0][0][2] [12]), 
      .C1(\buffer[12][0][2] [12]), .C2(n_27), .ZN(n_22_22_108));
   NAND4_X1 i_22_22_122 (.A1(n_22_22_115), .A2(n_22_22_113), .A3(n_22_22_111), 
      .A4(n_22_22_110), .ZN(n_22_22_109));
   AOI22_X1 i_22_22_123 (.A1(\buffer[15][0][2] [12]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][2] [12]), .ZN(n_22_22_110));
   AOI22_X1 i_22_22_124 (.A1(\buffer[10][0][2] [12]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][2] [12]), .ZN(n_22_22_111));
   AOI22_X1 i_22_22_125 (.A1(\buffer[6][0][2] [12]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][2] [12]), .ZN(n_22_22_112));
   AOI22_X1 i_22_22_126 (.A1(\buffer[9][0][2] [12]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][2] [12]), .ZN(n_22_22_113));
   AOI22_X1 i_22_22_127 (.A1(\buffer[14][0][2] [12]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][2] [12]), .ZN(n_22_22_114));
   AOI22_X1 i_22_22_128 (.A1(\buffer[11][0][2] [12]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][2] [12]), .ZN(n_22_22_115));
   AOI22_X1 i_22_22_129 (.A1(\buffer[13][0][2] [12]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][2] [12]), .ZN(n_22_22_116));
   NAND4_X1 i_22_22_130 (.A1(n_22_22_125), .A2(n_22_22_123), .A3(n_22_22_121), 
      .A4(n_22_22_117), .ZN(\output_filter[0][2] [13]));
   AOI221_X1 i_22_22_131 (.A(n_22_22_118), .B1(n_25), .B2(\buffer[0][0][2] [13]), 
      .C1(\buffer[12][0][2] [13]), .C2(n_27), .ZN(n_22_22_117));
   NAND4_X1 i_22_22_132 (.A1(n_22_22_124), .A2(n_22_22_122), .A3(n_22_22_120), 
      .A4(n_22_22_119), .ZN(n_22_22_118));
   AOI22_X1 i_22_22_133 (.A1(\buffer[15][0][2] [13]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][2] [13]), .ZN(n_22_22_119));
   AOI22_X1 i_22_22_134 (.A1(\buffer[10][0][2] [13]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][2] [13]), .ZN(n_22_22_120));
   AOI22_X1 i_22_22_135 (.A1(\buffer[6][0][2] [13]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][2] [13]), .ZN(n_22_22_121));
   AOI22_X1 i_22_22_136 (.A1(\buffer[9][0][2] [13]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][0][2] [13]), .ZN(n_22_22_122));
   AOI22_X1 i_22_22_137 (.A1(\buffer[14][0][2] [13]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][2] [13]), .ZN(n_22_22_123));
   AOI22_X1 i_22_22_138 (.A1(\buffer[11][0][2] [13]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][2] [13]), .ZN(n_22_22_124));
   AOI22_X1 i_22_22_139 (.A1(\buffer[13][0][2] [13]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][0][2] [13]), .ZN(n_22_22_125));
   NAND4_X1 i_22_22_140 (.A1(n_22_22_134), .A2(n_22_22_132), .A3(n_22_22_130), 
      .A4(n_22_22_126), .ZN(\output_filter[0][2] [14]));
   AOI221_X1 i_22_22_141 (.A(n_22_22_127), .B1(n_25), .B2(\buffer[0][0][2] [14]), 
      .C1(\buffer[12][0][2] [14]), .C2(n_27), .ZN(n_22_22_126));
   NAND4_X1 i_22_22_142 (.A1(n_22_22_133), .A2(n_22_22_131), .A3(n_22_22_129), 
      .A4(n_22_22_128), .ZN(n_22_22_127));
   AOI22_X1 i_22_22_143 (.A1(\buffer[15][0][2] [14]), .A2(n_22), .B1(n_16), 
      .B2(\buffer[8][0][2] [14]), .ZN(n_22_22_128));
   AOI22_X1 i_22_22_144 (.A1(\buffer[10][0][2] [14]), .A2(n_21), .B1(n_29), 
      .B2(\buffer[7][0][2] [14]), .ZN(n_22_22_129));
   AOI22_X1 i_22_22_145 (.A1(\buffer[6][0][2] [14]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][2] [14]), .ZN(n_22_22_130));
   AOI22_X1 i_22_22_146 (.A1(\buffer[9][0][2] [14]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][2] [14]), .ZN(n_22_22_131));
   AOI22_X1 i_22_22_147 (.A1(\buffer[14][0][2] [14]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][2] [14]), .ZN(n_22_22_132));
   AOI22_X1 i_22_22_148 (.A1(\buffer[11][0][2] [14]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][2] [14]), .ZN(n_22_22_133));
   AOI22_X1 i_22_22_149 (.A1(\buffer[13][0][2] [14]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][2] [14]), .ZN(n_22_22_134));
   NAND2_X1 i_22_22_150 (.A1(n_22_22_137), .A2(n_22_22_135), .ZN(
      \output_filter[0][2] [15]));
   AOI221_X1 i_22_22_151 (.A(n_22_22_136), .B1(n_31), .B2(\buffer[3][0][2] [15]), 
      .C1(\buffer[14][0][2] [15]), .C2(n_19), .ZN(n_22_22_135));
   NAND3_X1 i_22_22_152 (.A1(n_22_22_143), .A2(n_22_22_141), .A3(n_22_22_139), 
      .ZN(n_22_22_136));
   AOI221_X1 i_22_22_153 (.A(n_22_22_138), .B1(n_16), .B2(\buffer[8][0][2] [15]), 
      .C1(\buffer[13][0][2] [15]), .C2(n_26), .ZN(n_22_22_137));
   NAND3_X1 i_22_22_154 (.A1(n_22_22_144), .A2(n_22_22_142), .A3(n_22_22_140), 
      .ZN(n_22_22_138));
   AOI22_X1 i_22_22_155 (.A1(\buffer[11][0][2] [15]), .A2(n_17), .B1(n_24), 
      .B2(\buffer[2][0][2] [15]), .ZN(n_22_22_139));
   AOI22_X1 i_22_22_156 (.A1(\buffer[10][0][2] [15]), .A2(n_21), .B1(n_23), 
      .B2(\buffer[1][0][2] [15]), .ZN(n_22_22_140));
   AOI22_X1 i_22_22_157 (.A1(\buffer[6][0][2] [15]), .A2(n_28), .B1(n_18), 
      .B2(\buffer[5][0][2] [15]), .ZN(n_22_22_141));
   AOI22_X1 i_22_22_158 (.A1(\buffer[9][0][2] [15]), .A2(n_20), .B1(n_30), 
      .B2(\buffer[4][0][2] [15]), .ZN(n_22_22_142));
   AOI22_X1 i_22_22_159 (.A1(\buffer[7][0][2] [15]), .A2(n_29), .B1(n_25), 
      .B2(\buffer[0][0][2] [15]), .ZN(n_22_22_143));
   AOI22_X1 i_22_22_160 (.A1(\buffer[15][0][2] [15]), .A2(n_22), .B1(n_27), 
      .B2(\buffer[12][0][2] [15]), .ZN(n_22_22_144));
   NAND4_X1 i_21_21_0 (.A1(n_21_21_8), .A2(n_21_21_6), .A3(n_21_21_4), .A4(
      n_21_21_0), .ZN(\output_filter[0][1] [0]));
   AOI221_X1 i_21_21_1 (.A(n_21_21_1), .B1(n_25), .B2(\buffer[0][0][1] [0]), 
      .C1(\buffer[12][0][1] [0]), .C2(n_27), .ZN(n_21_21_0));
   NAND4_X1 i_21_21_2 (.A1(n_21_21_7), .A2(n_21_21_5), .A3(n_21_21_3), .A4(
      n_21_21_2), .ZN(n_21_21_1));
   AOI22_X1 i_21_21_3 (.A1(\buffer[15][0][1] [0]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][1] [0]), .ZN(n_21_21_2));
   AOI22_X1 i_21_21_4 (.A1(\buffer[10][0][1] [0]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][1] [0]), .ZN(n_21_21_3));
   AOI22_X1 i_21_21_5 (.A1(\buffer[6][0][1] [0]), .A2(n_28), .B1(n_30), .B2(
      \buffer[4][0][1] [0]), .ZN(n_21_21_4));
   AOI22_X1 i_21_21_6 (.A1(\buffer[9][0][1] [0]), .A2(n_20), .B1(n_31), .B2(
      \buffer[3][0][1] [0]), .ZN(n_21_21_5));
   AOI22_X1 i_21_21_7 (.A1(\buffer[14][0][1] [0]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][1] [0]), .ZN(n_21_21_6));
   AOI22_X1 i_21_21_8 (.A1(\buffer[11][0][1] [0]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][1] [0]), .ZN(n_21_21_7));
   AOI22_X1 i_21_21_9 (.A1(\buffer[13][0][1] [0]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][1] [0]), .ZN(n_21_21_8));
   NAND4_X1 i_21_21_10 (.A1(n_21_21_17), .A2(n_21_21_15), .A3(n_21_21_13), 
      .A4(n_21_21_9), .ZN(\output_filter[0][1] [1]));
   AOI221_X1 i_21_21_11 (.A(n_21_21_10), .B1(n_25), .B2(\buffer[0][0][1] [1]), 
      .C1(\buffer[12][0][1] [1]), .C2(n_27), .ZN(n_21_21_9));
   NAND4_X1 i_21_21_12 (.A1(n_21_21_16), .A2(n_21_21_14), .A3(n_21_21_12), 
      .A4(n_21_21_11), .ZN(n_21_21_10));
   AOI22_X1 i_21_21_13 (.A1(\buffer[15][0][1] [1]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][1] [1]), .ZN(n_21_21_11));
   AOI22_X1 i_21_21_14 (.A1(\buffer[10][0][1] [1]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][1] [1]), .ZN(n_21_21_12));
   AOI22_X1 i_21_21_15 (.A1(\buffer[6][0][1] [1]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][1] [1]), .ZN(n_21_21_13));
   AOI22_X1 i_21_21_16 (.A1(\buffer[9][0][1] [1]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][1] [1]), .ZN(n_21_21_14));
   AOI22_X1 i_21_21_17 (.A1(\buffer[14][0][1] [1]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][1] [1]), .ZN(n_21_21_15));
   AOI22_X1 i_21_21_18 (.A1(\buffer[11][0][1] [1]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][1] [1]), .ZN(n_21_21_16));
   AOI22_X1 i_21_21_19 (.A1(\buffer[13][0][1] [1]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][1] [1]), .ZN(n_21_21_17));
   NAND4_X1 i_21_21_20 (.A1(n_21_21_26), .A2(n_21_21_24), .A3(n_21_21_22), 
      .A4(n_21_21_18), .ZN(\output_filter[0][1] [2]));
   AOI221_X1 i_21_21_21 (.A(n_21_21_19), .B1(n_25), .B2(\buffer[0][0][1] [2]), 
      .C1(\buffer[12][0][1] [2]), .C2(n_27), .ZN(n_21_21_18));
   NAND4_X1 i_21_21_22 (.A1(n_21_21_25), .A2(n_21_21_23), .A3(n_21_21_21), 
      .A4(n_21_21_20), .ZN(n_21_21_19));
   AOI22_X1 i_21_21_23 (.A1(\buffer[15][0][1] [2]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][1] [2]), .ZN(n_21_21_20));
   AOI22_X1 i_21_21_24 (.A1(\buffer[10][0][1] [2]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][1] [2]), .ZN(n_21_21_21));
   AOI22_X1 i_21_21_25 (.A1(\buffer[6][0][1] [2]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][1] [2]), .ZN(n_21_21_22));
   AOI22_X1 i_21_21_26 (.A1(\buffer[9][0][1] [2]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][1] [2]), .ZN(n_21_21_23));
   AOI22_X1 i_21_21_27 (.A1(\buffer[14][0][1] [2]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][1] [2]), .ZN(n_21_21_24));
   AOI22_X1 i_21_21_28 (.A1(\buffer[11][0][1] [2]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][1] [2]), .ZN(n_21_21_25));
   AOI22_X1 i_21_21_29 (.A1(\buffer[13][0][1] [2]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][1] [2]), .ZN(n_21_21_26));
   NAND4_X1 i_21_21_30 (.A1(n_21_21_35), .A2(n_21_21_33), .A3(n_21_21_31), 
      .A4(n_21_21_27), .ZN(\output_filter[0][1] [3]));
   AOI221_X1 i_21_21_31 (.A(n_21_21_28), .B1(n_25), .B2(\buffer[0][0][1] [3]), 
      .C1(\buffer[12][0][1] [3]), .C2(n_27), .ZN(n_21_21_27));
   NAND4_X1 i_21_21_32 (.A1(n_21_21_34), .A2(n_21_21_32), .A3(n_21_21_30), 
      .A4(n_21_21_29), .ZN(n_21_21_28));
   AOI22_X1 i_21_21_33 (.A1(\buffer[15][0][1] [3]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][1] [3]), .ZN(n_21_21_29));
   AOI22_X1 i_21_21_34 (.A1(\buffer[10][0][1] [3]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][1] [3]), .ZN(n_21_21_30));
   AOI22_X1 i_21_21_35 (.A1(\buffer[6][0][1] [3]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][1] [3]), .ZN(n_21_21_31));
   AOI22_X1 i_21_21_36 (.A1(\buffer[9][0][1] [3]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][1] [3]), .ZN(n_21_21_32));
   AOI22_X1 i_21_21_37 (.A1(\buffer[14][0][1] [3]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][1] [3]), .ZN(n_21_21_33));
   AOI22_X1 i_21_21_38 (.A1(\buffer[11][0][1] [3]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][1] [3]), .ZN(n_21_21_34));
   AOI22_X1 i_21_21_39 (.A1(\buffer[13][0][1] [3]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][1] [3]), .ZN(n_21_21_35));
   NAND4_X1 i_21_21_40 (.A1(n_21_21_44), .A2(n_21_21_42), .A3(n_21_21_40), 
      .A4(n_21_21_36), .ZN(\output_filter[0][1] [4]));
   AOI221_X1 i_21_21_41 (.A(n_21_21_37), .B1(n_25), .B2(\buffer[0][0][1] [4]), 
      .C1(\buffer[12][0][1] [4]), .C2(n_27), .ZN(n_21_21_36));
   NAND4_X1 i_21_21_42 (.A1(n_21_21_43), .A2(n_21_21_41), .A3(n_21_21_39), 
      .A4(n_21_21_38), .ZN(n_21_21_37));
   AOI22_X1 i_21_21_43 (.A1(\buffer[15][0][1] [4]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][1] [4]), .ZN(n_21_21_38));
   AOI22_X1 i_21_21_44 (.A1(\buffer[10][0][1] [4]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][1] [4]), .ZN(n_21_21_39));
   AOI22_X1 i_21_21_45 (.A1(\buffer[6][0][1] [4]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][1] [4]), .ZN(n_21_21_40));
   AOI22_X1 i_21_21_46 (.A1(\buffer[9][0][1] [4]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][0][1] [4]), .ZN(n_21_21_41));
   AOI22_X1 i_21_21_47 (.A1(\buffer[14][0][1] [4]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][1] [4]), .ZN(n_21_21_42));
   AOI22_X1 i_21_21_48 (.A1(\buffer[11][0][1] [4]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][1] [4]), .ZN(n_21_21_43));
   AOI22_X1 i_21_21_49 (.A1(\buffer[13][0][1] [4]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][0][1] [4]), .ZN(n_21_21_44));
   NAND4_X1 i_21_21_50 (.A1(n_21_21_53), .A2(n_21_21_51), .A3(n_21_21_49), 
      .A4(n_21_21_45), .ZN(\output_filter[0][1] [5]));
   AOI221_X1 i_21_21_51 (.A(n_21_21_46), .B1(n_25), .B2(\buffer[0][0][1] [5]), 
      .C1(\buffer[12][0][1] [5]), .C2(n_27), .ZN(n_21_21_45));
   NAND4_X1 i_21_21_52 (.A1(n_21_21_52), .A2(n_21_21_50), .A3(n_21_21_48), 
      .A4(n_21_21_47), .ZN(n_21_21_46));
   AOI22_X1 i_21_21_53 (.A1(\buffer[15][0][1] [5]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][1] [5]), .ZN(n_21_21_47));
   AOI22_X1 i_21_21_54 (.A1(\buffer[10][0][1] [5]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][1] [5]), .ZN(n_21_21_48));
   AOI22_X1 i_21_21_55 (.A1(\buffer[6][0][1] [5]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][1] [5]), .ZN(n_21_21_49));
   AOI22_X1 i_21_21_56 (.A1(\buffer[9][0][1] [5]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][1] [5]), .ZN(n_21_21_50));
   AOI22_X1 i_21_21_57 (.A1(\buffer[14][0][1] [5]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][1] [5]), .ZN(n_21_21_51));
   AOI22_X1 i_21_21_58 (.A1(\buffer[11][0][1] [5]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][1] [5]), .ZN(n_21_21_52));
   AOI22_X1 i_21_21_59 (.A1(\buffer[13][0][1] [5]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][1] [5]), .ZN(n_21_21_53));
   NAND4_X1 i_21_21_60 (.A1(n_21_21_62), .A2(n_21_21_60), .A3(n_21_21_58), 
      .A4(n_21_21_54), .ZN(\output_filter[0][1] [6]));
   AOI221_X1 i_21_21_61 (.A(n_21_21_55), .B1(n_25), .B2(\buffer[0][0][1] [6]), 
      .C1(\buffer[12][0][1] [6]), .C2(n_27), .ZN(n_21_21_54));
   NAND4_X1 i_21_21_62 (.A1(n_21_21_61), .A2(n_21_21_59), .A3(n_21_21_57), 
      .A4(n_21_21_56), .ZN(n_21_21_55));
   AOI22_X1 i_21_21_63 (.A1(\buffer[15][0][1] [6]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][1] [6]), .ZN(n_21_21_56));
   AOI22_X1 i_21_21_64 (.A1(\buffer[10][0][1] [6]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][1] [6]), .ZN(n_21_21_57));
   AOI22_X1 i_21_21_65 (.A1(\buffer[6][0][1] [6]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][1] [6]), .ZN(n_21_21_58));
   AOI22_X1 i_21_21_66 (.A1(\buffer[9][0][1] [6]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][1] [6]), .ZN(n_21_21_59));
   AOI22_X1 i_21_21_67 (.A1(\buffer[14][0][1] [6]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][1] [6]), .ZN(n_21_21_60));
   AOI22_X1 i_21_21_68 (.A1(\buffer[11][0][1] [6]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][1] [6]), .ZN(n_21_21_61));
   AOI22_X1 i_21_21_69 (.A1(\buffer[13][0][1] [6]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][1] [6]), .ZN(n_21_21_62));
   NAND4_X1 i_21_21_70 (.A1(n_21_21_71), .A2(n_21_21_69), .A3(n_21_21_67), 
      .A4(n_21_21_63), .ZN(\output_filter[0][1] [7]));
   AOI221_X1 i_21_21_71 (.A(n_21_21_64), .B1(n_25), .B2(\buffer[0][0][1] [7]), 
      .C1(\buffer[12][0][1] [7]), .C2(n_27), .ZN(n_21_21_63));
   NAND4_X1 i_21_21_72 (.A1(n_21_21_70), .A2(n_21_21_68), .A3(n_21_21_66), 
      .A4(n_21_21_65), .ZN(n_21_21_64));
   AOI22_X1 i_21_21_73 (.A1(\buffer[15][0][1] [7]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][1] [7]), .ZN(n_21_21_65));
   AOI22_X1 i_21_21_74 (.A1(\buffer[10][0][1] [7]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][1] [7]), .ZN(n_21_21_66));
   AOI22_X1 i_21_21_75 (.A1(\buffer[6][0][1] [7]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][1] [7]), .ZN(n_21_21_67));
   AOI22_X1 i_21_21_76 (.A1(\buffer[9][0][1] [7]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][0][1] [7]), .ZN(n_21_21_68));
   AOI22_X1 i_21_21_77 (.A1(\buffer[14][0][1] [7]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][1] [7]), .ZN(n_21_21_69));
   AOI22_X1 i_21_21_78 (.A1(\buffer[11][0][1] [7]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][1] [7]), .ZN(n_21_21_70));
   AOI22_X1 i_21_21_79 (.A1(\buffer[13][0][1] [7]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][0][1] [7]), .ZN(n_21_21_71));
   NAND4_X1 i_21_21_80 (.A1(n_21_21_80), .A2(n_21_21_78), .A3(n_21_21_76), 
      .A4(n_21_21_72), .ZN(\output_filter[0][1] [8]));
   AOI221_X1 i_21_21_81 (.A(n_21_21_73), .B1(n_25), .B2(\buffer[0][0][1] [8]), 
      .C1(\buffer[12][0][1] [8]), .C2(n_27), .ZN(n_21_21_72));
   NAND4_X1 i_21_21_82 (.A1(n_21_21_79), .A2(n_21_21_77), .A3(n_21_21_75), 
      .A4(n_21_21_74), .ZN(n_21_21_73));
   AOI22_X1 i_21_21_83 (.A1(\buffer[15][0][1] [8]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][1] [8]), .ZN(n_21_21_74));
   AOI22_X1 i_21_21_84 (.A1(\buffer[10][0][1] [8]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][1] [8]), .ZN(n_21_21_75));
   AOI22_X1 i_21_21_85 (.A1(\buffer[6][0][1] [8]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][1] [8]), .ZN(n_21_21_76));
   AOI22_X1 i_21_21_86 (.A1(\buffer[9][0][1] [8]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][1] [8]), .ZN(n_21_21_77));
   AOI22_X1 i_21_21_87 (.A1(\buffer[14][0][1] [8]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][1] [8]), .ZN(n_21_21_78));
   AOI22_X1 i_21_21_88 (.A1(\buffer[11][0][1] [8]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][1] [8]), .ZN(n_21_21_79));
   AOI22_X1 i_21_21_89 (.A1(\buffer[13][0][1] [8]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][1] [8]), .ZN(n_21_21_80));
   NAND4_X1 i_21_21_90 (.A1(n_21_21_89), .A2(n_21_21_87), .A3(n_21_21_85), 
      .A4(n_21_21_81), .ZN(\output_filter[0][1] [9]));
   AOI221_X1 i_21_21_91 (.A(n_21_21_82), .B1(n_25), .B2(\buffer[0][0][1] [9]), 
      .C1(\buffer[12][0][1] [9]), .C2(n_27), .ZN(n_21_21_81));
   NAND4_X1 i_21_21_92 (.A1(n_21_21_88), .A2(n_21_21_86), .A3(n_21_21_84), 
      .A4(n_21_21_83), .ZN(n_21_21_82));
   AOI22_X1 i_21_21_93 (.A1(\buffer[15][0][1] [9]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][1] [9]), .ZN(n_21_21_83));
   AOI22_X1 i_21_21_94 (.A1(\buffer[10][0][1] [9]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][1] [9]), .ZN(n_21_21_84));
   AOI22_X1 i_21_21_95 (.A1(\buffer[6][0][1] [9]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][1] [9]), .ZN(n_21_21_85));
   AOI22_X1 i_21_21_96 (.A1(\buffer[9][0][1] [9]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][0][1] [9]), .ZN(n_21_21_86));
   AOI22_X1 i_21_21_97 (.A1(\buffer[14][0][1] [9]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][1] [9]), .ZN(n_21_21_87));
   AOI22_X1 i_21_21_98 (.A1(\buffer[11][0][1] [9]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][1] [9]), .ZN(n_21_21_88));
   AOI22_X1 i_21_21_99 (.A1(\buffer[13][0][1] [9]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][0][1] [9]), .ZN(n_21_21_89));
   NAND4_X1 i_21_21_100 (.A1(n_21_21_98), .A2(n_21_21_96), .A3(n_21_21_94), 
      .A4(n_21_21_90), .ZN(\output_filter[0][1] [10]));
   AOI221_X1 i_21_21_101 (.A(n_21_21_91), .B1(n_25), .B2(\buffer[0][0][1] [10]), 
      .C1(\buffer[12][0][1] [10]), .C2(n_27), .ZN(n_21_21_90));
   NAND4_X1 i_21_21_102 (.A1(n_21_21_97), .A2(n_21_21_95), .A3(n_21_21_93), 
      .A4(n_21_21_92), .ZN(n_21_21_91));
   AOI22_X1 i_21_21_103 (.A1(\buffer[15][0][1] [10]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][1] [10]), .ZN(n_21_21_92));
   AOI22_X1 i_21_21_104 (.A1(\buffer[10][0][1] [10]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][1] [10]), .ZN(n_21_21_93));
   AOI22_X1 i_21_21_105 (.A1(\buffer[6][0][1] [10]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][1] [10]), .ZN(n_21_21_94));
   AOI22_X1 i_21_21_106 (.A1(\buffer[9][0][1] [10]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][1] [10]), .ZN(n_21_21_95));
   AOI22_X1 i_21_21_107 (.A1(\buffer[14][0][1] [10]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][1] [10]), .ZN(n_21_21_96));
   AOI22_X1 i_21_21_108 (.A1(\buffer[11][0][1] [10]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][1] [10]), .ZN(n_21_21_97));
   AOI22_X1 i_21_21_109 (.A1(\buffer[13][0][1] [10]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][1] [10]), .ZN(n_21_21_98));
   NAND4_X1 i_21_21_110 (.A1(n_21_21_107), .A2(n_21_21_105), .A3(n_21_21_103), 
      .A4(n_21_21_99), .ZN(\output_filter[0][1] [11]));
   AOI221_X1 i_21_21_111 (.A(n_21_21_100), .B1(n_25), .B2(\buffer[0][0][1] [11]), 
      .C1(\buffer[12][0][1] [11]), .C2(n_27), .ZN(n_21_21_99));
   NAND4_X1 i_21_21_112 (.A1(n_21_21_106), .A2(n_21_21_104), .A3(n_21_21_102), 
      .A4(n_21_21_101), .ZN(n_21_21_100));
   AOI22_X1 i_21_21_113 (.A1(\buffer[15][0][1] [11]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][1] [11]), .ZN(n_21_21_101));
   AOI22_X1 i_21_21_114 (.A1(\buffer[10][0][1] [11]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][1] [11]), .ZN(n_21_21_102));
   AOI22_X1 i_21_21_115 (.A1(\buffer[6][0][1] [11]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][1] [11]), .ZN(n_21_21_103));
   AOI22_X1 i_21_21_116 (.A1(\buffer[9][0][1] [11]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][0][1] [11]), .ZN(n_21_21_104));
   AOI22_X1 i_21_21_117 (.A1(\buffer[14][0][1] [11]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][1] [11]), .ZN(n_21_21_105));
   AOI22_X1 i_21_21_118 (.A1(\buffer[11][0][1] [11]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][1] [11]), .ZN(n_21_21_106));
   AOI22_X1 i_21_21_119 (.A1(\buffer[13][0][1] [11]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][0][1] [11]), .ZN(n_21_21_107));
   NAND4_X1 i_21_21_120 (.A1(n_21_21_116), .A2(n_21_21_114), .A3(n_21_21_112), 
      .A4(n_21_21_108), .ZN(\output_filter[0][1] [12]));
   AOI221_X1 i_21_21_121 (.A(n_21_21_109), .B1(n_25), .B2(\buffer[0][0][1] [12]), 
      .C1(\buffer[12][0][1] [12]), .C2(n_27), .ZN(n_21_21_108));
   NAND4_X1 i_21_21_122 (.A1(n_21_21_115), .A2(n_21_21_113), .A3(n_21_21_111), 
      .A4(n_21_21_110), .ZN(n_21_21_109));
   AOI22_X1 i_21_21_123 (.A1(\buffer[15][0][1] [12]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][1] [12]), .ZN(n_21_21_110));
   AOI22_X1 i_21_21_124 (.A1(\buffer[10][0][1] [12]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][1] [12]), .ZN(n_21_21_111));
   AOI22_X1 i_21_21_125 (.A1(\buffer[6][0][1] [12]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][1] [12]), .ZN(n_21_21_112));
   AOI22_X1 i_21_21_126 (.A1(\buffer[9][0][1] [12]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][1] [12]), .ZN(n_21_21_113));
   AOI22_X1 i_21_21_127 (.A1(\buffer[14][0][1] [12]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][1] [12]), .ZN(n_21_21_114));
   AOI22_X1 i_21_21_128 (.A1(\buffer[11][0][1] [12]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][1] [12]), .ZN(n_21_21_115));
   AOI22_X1 i_21_21_129 (.A1(\buffer[13][0][1] [12]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][1] [12]), .ZN(n_21_21_116));
   NAND4_X1 i_21_21_130 (.A1(n_21_21_125), .A2(n_21_21_123), .A3(n_21_21_121), 
      .A4(n_21_21_117), .ZN(\output_filter[0][1] [13]));
   AOI221_X1 i_21_21_131 (.A(n_21_21_118), .B1(n_25), .B2(\buffer[0][0][1] [13]), 
      .C1(\buffer[12][0][1] [13]), .C2(n_27), .ZN(n_21_21_117));
   NAND4_X1 i_21_21_132 (.A1(n_21_21_124), .A2(n_21_21_122), .A3(n_21_21_120), 
      .A4(n_21_21_119), .ZN(n_21_21_118));
   AOI22_X1 i_21_21_133 (.A1(\buffer[15][0][1] [13]), .A2(n_22), .B1(n_29), 
      .B2(\buffer[7][0][1] [13]), .ZN(n_21_21_119));
   AOI22_X1 i_21_21_134 (.A1(\buffer[10][0][1] [13]), .A2(n_21), .B1(n_16), 
      .B2(\buffer[8][0][1] [13]), .ZN(n_21_21_120));
   AOI22_X1 i_21_21_135 (.A1(\buffer[6][0][1] [13]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][1] [13]), .ZN(n_21_21_121));
   AOI22_X1 i_21_21_136 (.A1(\buffer[9][0][1] [13]), .A2(n_20), .B1(n_24), 
      .B2(\buffer[2][0][1] [13]), .ZN(n_21_21_122));
   AOI22_X1 i_21_21_137 (.A1(\buffer[14][0][1] [13]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][1] [13]), .ZN(n_21_21_123));
   AOI22_X1 i_21_21_138 (.A1(\buffer[11][0][1] [13]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][1] [13]), .ZN(n_21_21_124));
   AOI22_X1 i_21_21_139 (.A1(\buffer[13][0][1] [13]), .A2(n_26), .B1(n_31), 
      .B2(\buffer[3][0][1] [13]), .ZN(n_21_21_125));
   NAND4_X1 i_21_21_140 (.A1(n_21_21_134), .A2(n_21_21_132), .A3(n_21_21_130), 
      .A4(n_21_21_126), .ZN(\output_filter[0][1] [14]));
   AOI221_X1 i_21_21_141 (.A(n_21_21_127), .B1(n_25), .B2(\buffer[0][0][1] [14]), 
      .C1(\buffer[12][0][1] [14]), .C2(n_27), .ZN(n_21_21_126));
   NAND4_X1 i_21_21_142 (.A1(n_21_21_133), .A2(n_21_21_131), .A3(n_21_21_129), 
      .A4(n_21_21_128), .ZN(n_21_21_127));
   AOI22_X1 i_21_21_143 (.A1(\buffer[15][0][1] [14]), .A2(n_22), .B1(n_16), 
      .B2(\buffer[8][0][1] [14]), .ZN(n_21_21_128));
   AOI22_X1 i_21_21_144 (.A1(\buffer[10][0][1] [14]), .A2(n_21), .B1(n_29), 
      .B2(\buffer[7][0][1] [14]), .ZN(n_21_21_129));
   AOI22_X1 i_21_21_145 (.A1(\buffer[6][0][1] [14]), .A2(n_28), .B1(n_30), 
      .B2(\buffer[4][0][1] [14]), .ZN(n_21_21_130));
   AOI22_X1 i_21_21_146 (.A1(\buffer[9][0][1] [14]), .A2(n_20), .B1(n_31), 
      .B2(\buffer[3][0][1] [14]), .ZN(n_21_21_131));
   AOI22_X1 i_21_21_147 (.A1(\buffer[14][0][1] [14]), .A2(n_19), .B1(n_23), 
      .B2(\buffer[1][0][1] [14]), .ZN(n_21_21_132));
   AOI22_X1 i_21_21_148 (.A1(\buffer[11][0][1] [14]), .A2(n_17), .B1(n_18), 
      .B2(\buffer[5][0][1] [14]), .ZN(n_21_21_133));
   AOI22_X1 i_21_21_149 (.A1(\buffer[13][0][1] [14]), .A2(n_26), .B1(n_24), 
      .B2(\buffer[2][0][1] [14]), .ZN(n_21_21_134));
   NAND2_X1 i_21_21_150 (.A1(n_21_21_137), .A2(n_21_21_135), .ZN(
      \output_filter[0][1] [15]));
   AOI221_X1 i_21_21_151 (.A(n_21_21_136), .B1(n_31), .B2(\buffer[3][0][1] [15]), 
      .C1(\buffer[14][0][1] [15]), .C2(n_19), .ZN(n_21_21_135));
   NAND3_X1 i_21_21_152 (.A1(n_21_21_143), .A2(n_21_21_141), .A3(n_21_21_139), 
      .ZN(n_21_21_136));
   AOI221_X1 i_21_21_153 (.A(n_21_21_138), .B1(n_16), .B2(\buffer[8][0][1] [15]), 
      .C1(\buffer[13][0][1] [15]), .C2(n_26), .ZN(n_21_21_137));
   NAND3_X1 i_21_21_154 (.A1(n_21_21_144), .A2(n_21_21_142), .A3(n_21_21_140), 
      .ZN(n_21_21_138));
   AOI22_X1 i_21_21_155 (.A1(\buffer[11][0][1] [15]), .A2(n_17), .B1(n_24), 
      .B2(\buffer[2][0][1] [15]), .ZN(n_21_21_139));
   AOI22_X1 i_21_21_156 (.A1(\buffer[10][0][1] [15]), .A2(n_21), .B1(n_23), 
      .B2(\buffer[1][0][1] [15]), .ZN(n_21_21_140));
   AOI22_X1 i_21_21_157 (.A1(\buffer[6][0][1] [15]), .A2(n_28), .B1(n_18), 
      .B2(\buffer[5][0][1] [15]), .ZN(n_21_21_141));
   AOI22_X1 i_21_21_158 (.A1(\buffer[9][0][1] [15]), .A2(n_20), .B1(n_30), 
      .B2(\buffer[4][0][1] [15]), .ZN(n_21_21_142));
   AOI22_X1 i_21_21_159 (.A1(\buffer[7][0][1] [15]), .A2(n_29), .B1(n_25), 
      .B2(\buffer[0][0][1] [15]), .ZN(n_21_21_143));
   AOI22_X1 i_21_21_160 (.A1(\buffer[15][0][1] [15]), .A2(n_22), .B1(n_27), 
      .B2(\buffer[12][0][1] [15]), .ZN(n_21_21_144));
   NAND2_X1 i_19_0_0 (.A1(n_19_0_2), .A2(n_19_0_0), .ZN(\output_filter[0][0] [0]));
   AOI221_X1 i_19_0_1 (.A(n_19_0_1), .B1(n_20), .B2(\buffer[9][0][0] [0]), 
      .C1(\buffer[10][0][0] [0]), .C2(n_21), .ZN(n_19_0_0));
   NAND3_X1 i_19_0_2 (.A1(n_19_0_8), .A2(n_19_0_6), .A3(n_19_0_4), .ZN(n_19_0_1));
   AOI221_X1 i_19_0_3 (.A(n_19_0_3), .B1(n_25), .B2(\buffer[0][0][0] [0]), 
      .C1(\buffer[2][0][0] [0]), .C2(n_24), .ZN(n_19_0_2));
   NAND3_X1 i_19_0_4 (.A1(n_19_0_9), .A2(n_19_0_7), .A3(n_19_0_5), .ZN(n_19_0_3));
   AOI22_X1 i_19_0_5 (.A1(\buffer[11][0][0] [0]), .A2(n_17), .B1(n_16), .B2(
      \buffer[8][0][0] [0]), .ZN(n_19_0_4));
   AOI22_X1 i_19_0_6 (.A1(\buffer[12][0][0] [0]), .A2(n_27), .B1(n_19), .B2(
      \buffer[14][0][0] [0]), .ZN(n_19_0_5));
   AOI22_X1 i_19_0_7 (.A1(\buffer[3][0][0] [0]), .A2(n_31), .B1(n_18), .B2(
      \buffer[5][0][0] [0]), .ZN(n_19_0_6));
   AOI22_X1 i_19_0_8 (.A1(\buffer[1][0][0] [0]), .A2(n_23), .B1(n_22), .B2(
      \buffer[15][0][0] [0]), .ZN(n_19_0_7));
   AOI22_X1 i_19_0_9 (.A1(\buffer[7][0][0] [0]), .A2(n_29), .B1(n_28), .B2(
      \buffer[6][0][0] [0]), .ZN(n_19_0_8));
   AOI22_X1 i_19_0_10 (.A1(\buffer[4][0][0] [0]), .A2(n_30), .B1(n_26), .B2(
      \buffer[13][0][0] [0]), .ZN(n_19_0_9));
   NAND2_X1 i_19_0_11 (.A1(n_19_0_12), .A2(n_19_0_10), .ZN(
      \output_filter[0][0] [1]));
   AOI221_X1 i_19_0_12 (.A(n_19_0_11), .B1(n_20), .B2(\buffer[9][0][0] [1]), 
      .C1(\buffer[10][0][0] [1]), .C2(n_21), .ZN(n_19_0_10));
   NAND3_X1 i_19_0_13 (.A1(n_19_0_18), .A2(n_19_0_16), .A3(n_19_0_14), .ZN(
      n_19_0_11));
   AOI221_X1 i_19_0_14 (.A(n_19_0_13), .B1(n_25), .B2(\buffer[0][0][0] [1]), 
      .C1(\buffer[2][0][0] [1]), .C2(n_24), .ZN(n_19_0_12));
   NAND3_X1 i_19_0_15 (.A1(n_19_0_19), .A2(n_19_0_17), .A3(n_19_0_15), .ZN(
      n_19_0_13));
   AOI22_X1 i_19_0_16 (.A1(\buffer[11][0][0] [1]), .A2(n_17), .B1(n_16), 
      .B2(\buffer[8][0][0] [1]), .ZN(n_19_0_14));
   AOI22_X1 i_19_0_17 (.A1(\buffer[12][0][0] [1]), .A2(n_27), .B1(n_19), 
      .B2(\buffer[14][0][0] [1]), .ZN(n_19_0_15));
   AOI22_X1 i_19_0_18 (.A1(\buffer[3][0][0] [1]), .A2(n_31), .B1(n_18), .B2(
      \buffer[5][0][0] [1]), .ZN(n_19_0_16));
   AOI22_X1 i_19_0_19 (.A1(\buffer[1][0][0] [1]), .A2(n_23), .B1(n_22), .B2(
      \buffer[15][0][0] [1]), .ZN(n_19_0_17));
   AOI22_X1 i_19_0_20 (.A1(\buffer[7][0][0] [1]), .A2(n_29), .B1(n_28), .B2(
      \buffer[6][0][0] [1]), .ZN(n_19_0_18));
   AOI22_X1 i_19_0_21 (.A1(\buffer[4][0][0] [1]), .A2(n_30), .B1(n_26), .B2(
      \buffer[13][0][0] [1]), .ZN(n_19_0_19));
   NAND2_X1 i_19_0_22 (.A1(n_19_0_22), .A2(n_19_0_20), .ZN(
      \output_filter[0][0] [2]));
   AOI221_X1 i_19_0_23 (.A(n_19_0_21), .B1(n_20), .B2(\buffer[9][0][0] [2]), 
      .C1(\buffer[10][0][0] [2]), .C2(n_21), .ZN(n_19_0_20));
   NAND3_X1 i_19_0_24 (.A1(n_19_0_28), .A2(n_19_0_26), .A3(n_19_0_24), .ZN(
      n_19_0_21));
   AOI221_X1 i_19_0_25 (.A(n_19_0_23), .B1(n_25), .B2(\buffer[0][0][0] [2]), 
      .C1(\buffer[2][0][0] [2]), .C2(n_24), .ZN(n_19_0_22));
   NAND3_X1 i_19_0_26 (.A1(n_19_0_29), .A2(n_19_0_27), .A3(n_19_0_25), .ZN(
      n_19_0_23));
   AOI22_X1 i_19_0_27 (.A1(\buffer[11][0][0] [2]), .A2(n_17), .B1(n_16), 
      .B2(\buffer[8][0][0] [2]), .ZN(n_19_0_24));
   AOI22_X1 i_19_0_28 (.A1(\buffer[12][0][0] [2]), .A2(n_27), .B1(n_19), 
      .B2(\buffer[14][0][0] [2]), .ZN(n_19_0_25));
   AOI22_X1 i_19_0_29 (.A1(\buffer[3][0][0] [2]), .A2(n_31), .B1(n_18), .B2(
      \buffer[5][0][0] [2]), .ZN(n_19_0_26));
   AOI22_X1 i_19_0_30 (.A1(\buffer[1][0][0] [2]), .A2(n_23), .B1(n_22), .B2(
      \buffer[15][0][0] [2]), .ZN(n_19_0_27));
   AOI22_X1 i_19_0_31 (.A1(\buffer[7][0][0] [2]), .A2(n_29), .B1(n_28), .B2(
      \buffer[6][0][0] [2]), .ZN(n_19_0_28));
   AOI22_X1 i_19_0_32 (.A1(\buffer[4][0][0] [2]), .A2(n_30), .B1(n_26), .B2(
      \buffer[13][0][0] [2]), .ZN(n_19_0_29));
   NAND2_X1 i_19_0_33 (.A1(n_19_0_32), .A2(n_19_0_30), .ZN(
      \output_filter[0][0] [3]));
   AOI221_X1 i_19_0_34 (.A(n_19_0_31), .B1(n_20), .B2(\buffer[9][0][0] [3]), 
      .C1(\buffer[10][0][0] [3]), .C2(n_21), .ZN(n_19_0_30));
   NAND3_X1 i_19_0_35 (.A1(n_19_0_38), .A2(n_19_0_36), .A3(n_19_0_34), .ZN(
      n_19_0_31));
   AOI221_X1 i_19_0_36 (.A(n_19_0_33), .B1(n_25), .B2(\buffer[0][0][0] [3]), 
      .C1(\buffer[2][0][0] [3]), .C2(n_24), .ZN(n_19_0_32));
   NAND3_X1 i_19_0_37 (.A1(n_19_0_39), .A2(n_19_0_37), .A3(n_19_0_35), .ZN(
      n_19_0_33));
   AOI22_X1 i_19_0_38 (.A1(\buffer[11][0][0] [3]), .A2(n_17), .B1(n_16), 
      .B2(\buffer[8][0][0] [3]), .ZN(n_19_0_34));
   AOI22_X1 i_19_0_39 (.A1(\buffer[12][0][0] [3]), .A2(n_27), .B1(n_19), 
      .B2(\buffer[14][0][0] [3]), .ZN(n_19_0_35));
   AOI22_X1 i_19_0_40 (.A1(\buffer[3][0][0] [3]), .A2(n_31), .B1(n_18), .B2(
      \buffer[5][0][0] [3]), .ZN(n_19_0_36));
   AOI22_X1 i_19_0_41 (.A1(\buffer[1][0][0] [3]), .A2(n_23), .B1(n_22), .B2(
      \buffer[15][0][0] [3]), .ZN(n_19_0_37));
   AOI22_X1 i_19_0_42 (.A1(\buffer[7][0][0] [3]), .A2(n_29), .B1(n_28), .B2(
      \buffer[6][0][0] [3]), .ZN(n_19_0_38));
   AOI22_X1 i_19_0_43 (.A1(\buffer[4][0][0] [3]), .A2(n_30), .B1(n_26), .B2(
      \buffer[13][0][0] [3]), .ZN(n_19_0_39));
   NAND2_X1 i_19_0_44 (.A1(n_19_0_42), .A2(n_19_0_40), .ZN(
      \output_filter[0][0] [4]));
   AOI221_X1 i_19_0_45 (.A(n_19_0_41), .B1(n_20), .B2(\buffer[9][0][0] [4]), 
      .C1(\buffer[10][0][0] [4]), .C2(n_21), .ZN(n_19_0_40));
   NAND3_X1 i_19_0_46 (.A1(n_19_0_48), .A2(n_19_0_46), .A3(n_19_0_44), .ZN(
      n_19_0_41));
   AOI221_X1 i_19_0_47 (.A(n_19_0_43), .B1(n_25), .B2(\buffer[0][0][0] [4]), 
      .C1(\buffer[3][0][0] [4]), .C2(n_31), .ZN(n_19_0_42));
   NAND3_X1 i_19_0_48 (.A1(n_19_0_49), .A2(n_19_0_47), .A3(n_19_0_45), .ZN(
      n_19_0_43));
   AOI22_X1 i_19_0_49 (.A1(\buffer[11][0][0] [4]), .A2(n_17), .B1(n_16), 
      .B2(\buffer[8][0][0] [4]), .ZN(n_19_0_44));
   AOI22_X1 i_19_0_50 (.A1(\buffer[12][0][0] [4]), .A2(n_27), .B1(n_19), 
      .B2(\buffer[14][0][0] [4]), .ZN(n_19_0_45));
   AOI22_X1 i_19_0_51 (.A1(\buffer[2][0][0] [4]), .A2(n_24), .B1(n_18), .B2(
      \buffer[5][0][0] [4]), .ZN(n_19_0_46));
   AOI22_X1 i_19_0_52 (.A1(\buffer[1][0][0] [4]), .A2(n_23), .B1(n_22), .B2(
      \buffer[15][0][0] [4]), .ZN(n_19_0_47));
   AOI22_X1 i_19_0_53 (.A1(\buffer[7][0][0] [4]), .A2(n_29), .B1(n_28), .B2(
      \buffer[6][0][0] [4]), .ZN(n_19_0_48));
   AOI22_X1 i_19_0_54 (.A1(\buffer[4][0][0] [4]), .A2(n_30), .B1(n_26), .B2(
      \buffer[13][0][0] [4]), .ZN(n_19_0_49));
   NAND2_X1 i_19_0_55 (.A1(n_19_0_52), .A2(n_19_0_50), .ZN(
      \output_filter[0][0] [5]));
   AOI221_X1 i_19_0_56 (.A(n_19_0_51), .B1(n_20), .B2(\buffer[9][0][0] [5]), 
      .C1(\buffer[10][0][0] [5]), .C2(n_21), .ZN(n_19_0_50));
   NAND3_X1 i_19_0_57 (.A1(n_19_0_58), .A2(n_19_0_56), .A3(n_19_0_54), .ZN(
      n_19_0_51));
   AOI221_X1 i_19_0_58 (.A(n_19_0_53), .B1(n_25), .B2(\buffer[0][0][0] [5]), 
      .C1(\buffer[2][0][0] [5]), .C2(n_24), .ZN(n_19_0_52));
   NAND3_X1 i_19_0_59 (.A1(n_19_0_59), .A2(n_19_0_57), .A3(n_19_0_55), .ZN(
      n_19_0_53));
   AOI22_X1 i_19_0_60 (.A1(\buffer[11][0][0] [5]), .A2(n_17), .B1(n_16), 
      .B2(\buffer[8][0][0] [5]), .ZN(n_19_0_54));
   AOI22_X1 i_19_0_61 (.A1(\buffer[12][0][0] [5]), .A2(n_27), .B1(n_19), 
      .B2(\buffer[14][0][0] [5]), .ZN(n_19_0_55));
   AOI22_X1 i_19_0_62 (.A1(\buffer[3][0][0] [5]), .A2(n_31), .B1(n_18), .B2(
      \buffer[5][0][0] [5]), .ZN(n_19_0_56));
   AOI22_X1 i_19_0_63 (.A1(\buffer[1][0][0] [5]), .A2(n_23), .B1(n_22), .B2(
      \buffer[15][0][0] [5]), .ZN(n_19_0_57));
   AOI22_X1 i_19_0_64 (.A1(\buffer[7][0][0] [5]), .A2(n_29), .B1(n_28), .B2(
      \buffer[6][0][0] [5]), .ZN(n_19_0_58));
   AOI22_X1 i_19_0_65 (.A1(\buffer[4][0][0] [5]), .A2(n_30), .B1(n_26), .B2(
      \buffer[13][0][0] [5]), .ZN(n_19_0_59));
   NAND2_X1 i_19_0_66 (.A1(n_19_0_62), .A2(n_19_0_60), .ZN(
      \output_filter[0][0] [6]));
   AOI221_X1 i_19_0_67 (.A(n_19_0_61), .B1(n_20), .B2(\buffer[9][0][0] [6]), 
      .C1(\buffer[10][0][0] [6]), .C2(n_21), .ZN(n_19_0_60));
   NAND3_X1 i_19_0_68 (.A1(n_19_0_68), .A2(n_19_0_66), .A3(n_19_0_64), .ZN(
      n_19_0_61));
   AOI221_X1 i_19_0_69 (.A(n_19_0_63), .B1(n_25), .B2(\buffer[0][0][0] [6]), 
      .C1(\buffer[2][0][0] [6]), .C2(n_24), .ZN(n_19_0_62));
   NAND3_X1 i_19_0_70 (.A1(n_19_0_69), .A2(n_19_0_67), .A3(n_19_0_65), .ZN(
      n_19_0_63));
   AOI22_X1 i_19_0_71 (.A1(\buffer[11][0][0] [6]), .A2(n_17), .B1(n_16), 
      .B2(\buffer[8][0][0] [6]), .ZN(n_19_0_64));
   AOI22_X1 i_19_0_72 (.A1(\buffer[12][0][0] [6]), .A2(n_27), .B1(n_19), 
      .B2(\buffer[14][0][0] [6]), .ZN(n_19_0_65));
   AOI22_X1 i_19_0_73 (.A1(\buffer[3][0][0] [6]), .A2(n_31), .B1(n_18), .B2(
      \buffer[5][0][0] [6]), .ZN(n_19_0_66));
   AOI22_X1 i_19_0_74 (.A1(\buffer[1][0][0] [6]), .A2(n_23), .B1(n_22), .B2(
      \buffer[15][0][0] [6]), .ZN(n_19_0_67));
   AOI22_X1 i_19_0_75 (.A1(\buffer[7][0][0] [6]), .A2(n_29), .B1(n_28), .B2(
      \buffer[6][0][0] [6]), .ZN(n_19_0_68));
   AOI22_X1 i_19_0_76 (.A1(\buffer[4][0][0] [6]), .A2(n_30), .B1(n_26), .B2(
      \buffer[13][0][0] [6]), .ZN(n_19_0_69));
   NAND2_X1 i_19_0_77 (.A1(n_19_0_72), .A2(n_19_0_70), .ZN(
      \output_filter[0][0] [7]));
   AOI221_X1 i_19_0_78 (.A(n_19_0_71), .B1(n_20), .B2(\buffer[9][0][0] [7]), 
      .C1(\buffer[10][0][0] [7]), .C2(n_21), .ZN(n_19_0_70));
   NAND3_X1 i_19_0_79 (.A1(n_19_0_78), .A2(n_19_0_76), .A3(n_19_0_74), .ZN(
      n_19_0_71));
   AOI221_X1 i_19_0_80 (.A(n_19_0_73), .B1(n_25), .B2(\buffer[0][0][0] [7]), 
      .C1(\buffer[3][0][0] [7]), .C2(n_31), .ZN(n_19_0_72));
   NAND3_X1 i_19_0_81 (.A1(n_19_0_79), .A2(n_19_0_77), .A3(n_19_0_75), .ZN(
      n_19_0_73));
   AOI22_X1 i_19_0_82 (.A1(\buffer[11][0][0] [7]), .A2(n_17), .B1(n_16), 
      .B2(\buffer[8][0][0] [7]), .ZN(n_19_0_74));
   AOI22_X1 i_19_0_83 (.A1(\buffer[12][0][0] [7]), .A2(n_27), .B1(n_19), 
      .B2(\buffer[14][0][0] [7]), .ZN(n_19_0_75));
   AOI22_X1 i_19_0_84 (.A1(\buffer[2][0][0] [7]), .A2(n_24), .B1(n_18), .B2(
      \buffer[5][0][0] [7]), .ZN(n_19_0_76));
   AOI22_X1 i_19_0_85 (.A1(\buffer[1][0][0] [7]), .A2(n_23), .B1(n_22), .B2(
      \buffer[15][0][0] [7]), .ZN(n_19_0_77));
   AOI22_X1 i_19_0_86 (.A1(\buffer[7][0][0] [7]), .A2(n_29), .B1(n_28), .B2(
      \buffer[6][0][0] [7]), .ZN(n_19_0_78));
   AOI22_X1 i_19_0_87 (.A1(\buffer[4][0][0] [7]), .A2(n_30), .B1(n_26), .B2(
      \buffer[13][0][0] [7]), .ZN(n_19_0_79));
   NAND2_X1 i_19_0_88 (.A1(n_19_0_82), .A2(n_19_0_80), .ZN(
      \output_filter[0][0] [8]));
   AOI221_X1 i_19_0_89 (.A(n_19_0_81), .B1(n_20), .B2(\buffer[9][0][0] [8]), 
      .C1(\buffer[10][0][0] [8]), .C2(n_21), .ZN(n_19_0_80));
   NAND3_X1 i_19_0_90 (.A1(n_19_0_88), .A2(n_19_0_86), .A3(n_19_0_84), .ZN(
      n_19_0_81));
   AOI221_X1 i_19_0_91 (.A(n_19_0_83), .B1(n_25), .B2(\buffer[0][0][0] [8]), 
      .C1(\buffer[2][0][0] [8]), .C2(n_24), .ZN(n_19_0_82));
   NAND3_X1 i_19_0_92 (.A1(n_19_0_89), .A2(n_19_0_87), .A3(n_19_0_85), .ZN(
      n_19_0_83));
   AOI22_X1 i_19_0_93 (.A1(\buffer[11][0][0] [8]), .A2(n_17), .B1(n_16), 
      .B2(\buffer[8][0][0] [8]), .ZN(n_19_0_84));
   AOI22_X1 i_19_0_94 (.A1(\buffer[12][0][0] [8]), .A2(n_27), .B1(n_19), 
      .B2(\buffer[14][0][0] [8]), .ZN(n_19_0_85));
   AOI22_X1 i_19_0_95 (.A1(\buffer[3][0][0] [8]), .A2(n_31), .B1(n_18), .B2(
      \buffer[5][0][0] [8]), .ZN(n_19_0_86));
   AOI22_X1 i_19_0_96 (.A1(\buffer[1][0][0] [8]), .A2(n_23), .B1(n_22), .B2(
      \buffer[15][0][0] [8]), .ZN(n_19_0_87));
   AOI22_X1 i_19_0_97 (.A1(\buffer[7][0][0] [8]), .A2(n_29), .B1(n_28), .B2(
      \buffer[6][0][0] [8]), .ZN(n_19_0_88));
   AOI22_X1 i_19_0_98 (.A1(\buffer[4][0][0] [8]), .A2(n_30), .B1(n_26), .B2(
      \buffer[13][0][0] [8]), .ZN(n_19_0_89));
   NAND2_X1 i_19_0_99 (.A1(n_19_0_92), .A2(n_19_0_90), .ZN(
      \output_filter[0][0] [9]));
   AOI221_X1 i_19_0_100 (.A(n_19_0_91), .B1(n_20), .B2(\buffer[9][0][0] [9]), 
      .C1(\buffer[10][0][0] [9]), .C2(n_21), .ZN(n_19_0_90));
   NAND3_X1 i_19_0_101 (.A1(n_19_0_98), .A2(n_19_0_96), .A3(n_19_0_94), .ZN(
      n_19_0_91));
   AOI221_X1 i_19_0_102 (.A(n_19_0_93), .B1(n_25), .B2(\buffer[0][0][0] [9]), 
      .C1(\buffer[3][0][0] [9]), .C2(n_31), .ZN(n_19_0_92));
   NAND3_X1 i_19_0_103 (.A1(n_19_0_99), .A2(n_19_0_97), .A3(n_19_0_95), .ZN(
      n_19_0_93));
   AOI22_X1 i_19_0_104 (.A1(\buffer[11][0][0] [9]), .A2(n_17), .B1(n_16), 
      .B2(\buffer[8][0][0] [9]), .ZN(n_19_0_94));
   AOI22_X1 i_19_0_105 (.A1(\buffer[12][0][0] [9]), .A2(n_27), .B1(n_19), 
      .B2(\buffer[14][0][0] [9]), .ZN(n_19_0_95));
   AOI22_X1 i_19_0_106 (.A1(\buffer[2][0][0] [9]), .A2(n_24), .B1(n_18), 
      .B2(\buffer[5][0][0] [9]), .ZN(n_19_0_96));
   AOI22_X1 i_19_0_107 (.A1(\buffer[1][0][0] [9]), .A2(n_23), .B1(n_22), 
      .B2(\buffer[15][0][0] [9]), .ZN(n_19_0_97));
   AOI22_X1 i_19_0_108 (.A1(\buffer[7][0][0] [9]), .A2(n_29), .B1(n_28), 
      .B2(\buffer[6][0][0] [9]), .ZN(n_19_0_98));
   AOI22_X1 i_19_0_109 (.A1(\buffer[4][0][0] [9]), .A2(n_30), .B1(n_26), 
      .B2(\buffer[13][0][0] [9]), .ZN(n_19_0_99));
   NAND2_X1 i_19_0_110 (.A1(n_19_0_102), .A2(n_19_0_100), .ZN(
      \output_filter[0][0] [10]));
   AOI221_X1 i_19_0_111 (.A(n_19_0_101), .B1(n_20), .B2(\buffer[9][0][0] [10]), 
      .C1(\buffer[10][0][0] [10]), .C2(n_21), .ZN(n_19_0_100));
   NAND3_X1 i_19_0_112 (.A1(n_19_0_108), .A2(n_19_0_106), .A3(n_19_0_104), 
      .ZN(n_19_0_101));
   AOI221_X1 i_19_0_113 (.A(n_19_0_103), .B1(n_25), .B2(\buffer[0][0][0] [10]), 
      .C1(\buffer[2][0][0] [10]), .C2(n_24), .ZN(n_19_0_102));
   NAND3_X1 i_19_0_114 (.A1(n_19_0_109), .A2(n_19_0_107), .A3(n_19_0_105), 
      .ZN(n_19_0_103));
   AOI22_X1 i_19_0_115 (.A1(\buffer[11][0][0] [10]), .A2(n_17), .B1(n_16), 
      .B2(\buffer[8][0][0] [10]), .ZN(n_19_0_104));
   AOI22_X1 i_19_0_116 (.A1(\buffer[12][0][0] [10]), .A2(n_27), .B1(n_19), 
      .B2(\buffer[14][0][0] [10]), .ZN(n_19_0_105));
   AOI22_X1 i_19_0_117 (.A1(\buffer[3][0][0] [10]), .A2(n_31), .B1(n_18), 
      .B2(\buffer[5][0][0] [10]), .ZN(n_19_0_106));
   AOI22_X1 i_19_0_118 (.A1(\buffer[1][0][0] [10]), .A2(n_23), .B1(n_22), 
      .B2(\buffer[15][0][0] [10]), .ZN(n_19_0_107));
   AOI22_X1 i_19_0_119 (.A1(\buffer[7][0][0] [10]), .A2(n_29), .B1(n_28), 
      .B2(\buffer[6][0][0] [10]), .ZN(n_19_0_108));
   AOI22_X1 i_19_0_120 (.A1(\buffer[4][0][0] [10]), .A2(n_30), .B1(n_26), 
      .B2(\buffer[13][0][0] [10]), .ZN(n_19_0_109));
   NAND2_X1 i_19_0_121 (.A1(n_19_0_112), .A2(n_19_0_110), .ZN(
      \output_filter[0][0] [11]));
   AOI221_X1 i_19_0_122 (.A(n_19_0_111), .B1(n_20), .B2(\buffer[9][0][0] [11]), 
      .C1(\buffer[10][0][0] [11]), .C2(n_21), .ZN(n_19_0_110));
   NAND3_X1 i_19_0_123 (.A1(n_19_0_118), .A2(n_19_0_116), .A3(n_19_0_114), 
      .ZN(n_19_0_111));
   AOI221_X1 i_19_0_124 (.A(n_19_0_113), .B1(n_25), .B2(\buffer[0][0][0] [11]), 
      .C1(\buffer[3][0][0] [11]), .C2(n_31), .ZN(n_19_0_112));
   NAND3_X1 i_19_0_125 (.A1(n_19_0_119), .A2(n_19_0_117), .A3(n_19_0_115), 
      .ZN(n_19_0_113));
   AOI22_X1 i_19_0_126 (.A1(\buffer[11][0][0] [11]), .A2(n_17), .B1(n_16), 
      .B2(\buffer[8][0][0] [11]), .ZN(n_19_0_114));
   AOI22_X1 i_19_0_127 (.A1(\buffer[12][0][0] [11]), .A2(n_27), .B1(n_19), 
      .B2(\buffer[14][0][0] [11]), .ZN(n_19_0_115));
   AOI22_X1 i_19_0_128 (.A1(\buffer[2][0][0] [11]), .A2(n_24), .B1(n_18), 
      .B2(\buffer[5][0][0] [11]), .ZN(n_19_0_116));
   AOI22_X1 i_19_0_129 (.A1(\buffer[1][0][0] [11]), .A2(n_23), .B1(n_22), 
      .B2(\buffer[15][0][0] [11]), .ZN(n_19_0_117));
   AOI22_X1 i_19_0_130 (.A1(\buffer[7][0][0] [11]), .A2(n_29), .B1(n_28), 
      .B2(\buffer[6][0][0] [11]), .ZN(n_19_0_118));
   AOI22_X1 i_19_0_131 (.A1(\buffer[4][0][0] [11]), .A2(n_30), .B1(n_26), 
      .B2(\buffer[13][0][0] [11]), .ZN(n_19_0_119));
   NAND2_X1 i_19_0_132 (.A1(n_19_0_122), .A2(n_19_0_120), .ZN(
      \output_filter[0][0] [12]));
   AOI221_X1 i_19_0_133 (.A(n_19_0_121), .B1(n_20), .B2(\buffer[9][0][0] [12]), 
      .C1(\buffer[10][0][0] [12]), .C2(n_21), .ZN(n_19_0_120));
   NAND3_X1 i_19_0_134 (.A1(n_19_0_128), .A2(n_19_0_126), .A3(n_19_0_124), 
      .ZN(n_19_0_121));
   AOI221_X1 i_19_0_135 (.A(n_19_0_123), .B1(n_25), .B2(\buffer[0][0][0] [12]), 
      .C1(\buffer[2][0][0] [12]), .C2(n_24), .ZN(n_19_0_122));
   NAND3_X1 i_19_0_136 (.A1(n_19_0_129), .A2(n_19_0_127), .A3(n_19_0_125), 
      .ZN(n_19_0_123));
   AOI22_X1 i_19_0_137 (.A1(\buffer[11][0][0] [12]), .A2(n_17), .B1(n_16), 
      .B2(\buffer[8][0][0] [12]), .ZN(n_19_0_124));
   AOI22_X1 i_19_0_138 (.A1(\buffer[12][0][0] [12]), .A2(n_27), .B1(n_19), 
      .B2(\buffer[14][0][0] [12]), .ZN(n_19_0_125));
   AOI22_X1 i_19_0_139 (.A1(\buffer[3][0][0] [12]), .A2(n_31), .B1(n_18), 
      .B2(\buffer[5][0][0] [12]), .ZN(n_19_0_126));
   AOI22_X1 i_19_0_140 (.A1(\buffer[1][0][0] [12]), .A2(n_23), .B1(n_22), 
      .B2(\buffer[15][0][0] [12]), .ZN(n_19_0_127));
   AOI22_X1 i_19_0_141 (.A1(\buffer[7][0][0] [12]), .A2(n_29), .B1(n_28), 
      .B2(\buffer[6][0][0] [12]), .ZN(n_19_0_128));
   AOI22_X1 i_19_0_142 (.A1(\buffer[4][0][0] [12]), .A2(n_30), .B1(n_26), 
      .B2(\buffer[13][0][0] [12]), .ZN(n_19_0_129));
   NAND2_X1 i_19_0_143 (.A1(n_19_0_132), .A2(n_19_0_130), .ZN(
      \output_filter[0][0] [13]));
   AOI221_X1 i_19_0_144 (.A(n_19_0_131), .B1(n_20), .B2(\buffer[9][0][0] [13]), 
      .C1(\buffer[10][0][0] [13]), .C2(n_21), .ZN(n_19_0_130));
   NAND3_X1 i_19_0_145 (.A1(n_19_0_138), .A2(n_19_0_136), .A3(n_19_0_134), 
      .ZN(n_19_0_131));
   AOI221_X1 i_19_0_146 (.A(n_19_0_133), .B1(n_25), .B2(\buffer[0][0][0] [13]), 
      .C1(\buffer[3][0][0] [13]), .C2(n_31), .ZN(n_19_0_132));
   NAND3_X1 i_19_0_147 (.A1(n_19_0_139), .A2(n_19_0_137), .A3(n_19_0_135), 
      .ZN(n_19_0_133));
   AOI22_X1 i_19_0_148 (.A1(\buffer[11][0][0] [13]), .A2(n_17), .B1(n_16), 
      .B2(\buffer[8][0][0] [13]), .ZN(n_19_0_134));
   AOI22_X1 i_19_0_149 (.A1(\buffer[12][0][0] [13]), .A2(n_27), .B1(n_19), 
      .B2(\buffer[14][0][0] [13]), .ZN(n_19_0_135));
   AOI22_X1 i_19_0_150 (.A1(\buffer[2][0][0] [13]), .A2(n_24), .B1(n_18), 
      .B2(\buffer[5][0][0] [13]), .ZN(n_19_0_136));
   AOI22_X1 i_19_0_151 (.A1(\buffer[1][0][0] [13]), .A2(n_23), .B1(n_22), 
      .B2(\buffer[15][0][0] [13]), .ZN(n_19_0_137));
   AOI22_X1 i_19_0_152 (.A1(\buffer[7][0][0] [13]), .A2(n_29), .B1(n_28), 
      .B2(\buffer[6][0][0] [13]), .ZN(n_19_0_138));
   AOI22_X1 i_19_0_153 (.A1(\buffer[4][0][0] [13]), .A2(n_30), .B1(n_26), 
      .B2(\buffer[13][0][0] [13]), .ZN(n_19_0_139));
   NAND2_X1 i_19_0_154 (.A1(n_19_0_142), .A2(n_19_0_140), .ZN(
      \output_filter[0][0] [14]));
   AOI221_X1 i_19_0_155 (.A(n_19_0_141), .B1(n_29), .B2(\buffer[7][0][0] [14]), 
      .C1(\buffer[10][0][0] [14]), .C2(n_21), .ZN(n_19_0_140));
   NAND3_X1 i_19_0_156 (.A1(n_19_0_148), .A2(n_19_0_146), .A3(n_19_0_144), 
      .ZN(n_19_0_141));
   AOI221_X1 i_19_0_157 (.A(n_19_0_143), .B1(n_25), .B2(\buffer[0][0][0] [14]), 
      .C1(\buffer[2][0][0] [14]), .C2(n_24), .ZN(n_19_0_142));
   NAND3_X1 i_19_0_158 (.A1(n_19_0_149), .A2(n_19_0_147), .A3(n_19_0_145), 
      .ZN(n_19_0_143));
   AOI22_X1 i_19_0_159 (.A1(\buffer[9][0][0] [14]), .A2(n_20), .B1(n_17), 
      .B2(\buffer[11][0][0] [14]), .ZN(n_19_0_144));
   AOI22_X1 i_19_0_160 (.A1(\buffer[12][0][0] [14]), .A2(n_27), .B1(n_19), 
      .B2(\buffer[14][0][0] [14]), .ZN(n_19_0_145));
   AOI22_X1 i_19_0_161 (.A1(\buffer[3][0][0] [14]), .A2(n_31), .B1(n_18), 
      .B2(\buffer[5][0][0] [14]), .ZN(n_19_0_146));
   AOI22_X1 i_19_0_162 (.A1(\buffer[1][0][0] [14]), .A2(n_23), .B1(n_22), 
      .B2(\buffer[15][0][0] [14]), .ZN(n_19_0_147));
   AOI22_X1 i_19_0_163 (.A1(\buffer[6][0][0] [14]), .A2(n_28), .B1(n_16), 
      .B2(\buffer[8][0][0] [14]), .ZN(n_19_0_148));
   AOI22_X1 i_19_0_164 (.A1(\buffer[4][0][0] [14]), .A2(n_30), .B1(n_26), 
      .B2(\buffer[13][0][0] [14]), .ZN(n_19_0_149));
   NAND2_X1 i_19_0_165 (.A1(n_19_0_152), .A2(n_19_0_150), .ZN(
      \output_filter[0][0] [15]));
   AOI221_X1 i_19_0_166 (.A(n_19_0_151), .B1(n_20), .B2(\buffer[9][0][0] [15]), 
      .C1(\buffer[10][0][0] [15]), .C2(n_21), .ZN(n_19_0_150));
   NAND3_X1 i_19_0_167 (.A1(n_19_0_161), .A2(n_19_0_157), .A3(n_19_0_154), 
      .ZN(n_19_0_151));
   AOI221_X1 i_19_0_168 (.A(n_19_0_153), .B1(n_18), .B2(\buffer[5][0][0] [15]), 
      .C1(\buffer[14][0][0] [15]), .C2(n_19), .ZN(n_19_0_152));
   NAND3_X1 i_19_0_169 (.A1(n_19_0_163), .A2(n_19_0_158), .A3(n_19_0_156), 
      .ZN(n_19_0_153));
   AOI22_X1 i_19_0_170 (.A1(\buffer[11][0][0] [15]), .A2(n_17), .B1(n_16), 
      .B2(\buffer[8][0][0] [15]), .ZN(n_19_0_154));
   NOR3_X1 i_19_0_171 (.A1(n_19_0_155), .A2(index_buffer[0]), .A3(
      index_buffer[1]), .ZN(n_16));
   NOR2_X1 i_19_0_172 (.A1(n_19_0_165), .A2(n_19_0_155), .ZN(n_17));
   NOR2_X1 i_19_0_173 (.A1(n_19_0_164), .A2(n_19_0_159), .ZN(n_18));
   NOR2_X1 i_19_0_174 (.A1(n_19_0_162), .A2(n_19_0_160), .ZN(n_19));
   NOR2_X1 i_19_0_175 (.A1(n_19_0_159), .A2(n_19_0_155), .ZN(n_20));
   NOR2_X1 i_19_0_176 (.A1(n_19_0_162), .A2(n_19_0_155), .ZN(n_21));
   OR2_X1 i_19_0_177 (.A1(n_19_0_167), .A2(index_buffer[2]), .ZN(n_19_0_155));
   AOI22_X1 i_19_0_178 (.A1(\buffer[1][0][0] [15]), .A2(n_23), .B1(n_22), 
      .B2(\buffer[15][0][0] [15]), .ZN(n_19_0_156));
   NOR2_X1 i_19_0_179 (.A1(n_19_0_165), .A2(n_19_0_160), .ZN(n_22));
   NOR3_X1 i_19_0_180 (.A1(n_19_0_159), .A2(index_buffer[2]), .A3(
      index_buffer[3]), .ZN(n_23));
   AOI22_X1 i_19_0_181 (.A1(\buffer[0][0][0] [15]), .A2(n_25), .B1(n_24), 
      .B2(\buffer[2][0][0] [15]), .ZN(n_19_0_157));
   NOR3_X1 i_19_0_182 (.A1(n_19_0_162), .A2(index_buffer[2]), .A3(
      index_buffer[3]), .ZN(n_24));
   NOR4_X1 i_19_0_183 (.A1(index_buffer[3]), .A2(index_buffer[2]), .A3(
      index_buffer[1]), .A4(index_buffer[0]), .ZN(n_25));
   AOI22_X1 i_19_0_184 (.A1(\buffer[12][0][0] [15]), .A2(n_27), .B1(n_26), 
      .B2(\buffer[13][0][0] [15]), .ZN(n_19_0_158));
   NOR2_X1 i_19_0_185 (.A1(n_19_0_160), .A2(n_19_0_159), .ZN(n_26));
   OR2_X1 i_19_0_186 (.A1(n_19_0_166), .A2(index_buffer[1]), .ZN(n_19_0_159));
   NOR3_X1 i_19_0_187 (.A1(n_19_0_160), .A2(index_buffer[0]), .A3(
      index_buffer[1]), .ZN(n_27));
   NAND2_X1 i_19_0_188 (.A1(index_buffer[3]), .A2(index_buffer[2]), .ZN(
      n_19_0_160));
   AOI22_X1 i_19_0_189 (.A1(\buffer[7][0][0] [15]), .A2(n_29), .B1(n_28), 
      .B2(\buffer[6][0][0] [15]), .ZN(n_19_0_161));
   NOR2_X1 i_19_0_190 (.A1(n_19_0_164), .A2(n_19_0_162), .ZN(n_28));
   NAND2_X1 i_19_0_191 (.A1(n_19_0_166), .A2(index_buffer[1]), .ZN(n_19_0_162));
   NOR2_X1 i_19_0_192 (.A1(n_19_0_165), .A2(n_19_0_164), .ZN(n_29));
   AOI22_X1 i_19_0_193 (.A1(\buffer[3][0][0] [15]), .A2(n_31), .B1(n_30), 
      .B2(\buffer[4][0][0] [15]), .ZN(n_19_0_163));
   NOR3_X1 i_19_0_194 (.A1(n_19_0_164), .A2(index_buffer[0]), .A3(
      index_buffer[1]), .ZN(n_30));
   NAND2_X1 i_19_0_195 (.A1(n_19_0_167), .A2(index_buffer[2]), .ZN(n_19_0_164));
   NOR3_X1 i_19_0_196 (.A1(n_19_0_165), .A2(index_buffer[2]), .A3(
      index_buffer[3]), .ZN(n_31));
   NAND2_X1 i_19_0_197 (.A1(index_buffer[1]), .A2(index_buffer[0]), .ZN(
      n_19_0_165));
   INV_X1 i_19_0_198 (.A(index_buffer[0]), .ZN(n_19_0_166));
   INV_X1 i_19_0_199 (.A(index_buffer[3]), .ZN(n_19_0_167));
endmodule

/* blackbox module Booth_Multiplier_bbox_23 */

/* blackbox module Booth_Multiplier_bbox_22 */

/* blackbox module Booth_Multiplier_bbox_21 */

/* blackbox module Booth_Multiplier_bbox_20 */

/* blackbox module Booth_Multiplier_bbox_19 */

/* blackbox module Booth_Multiplier_bbox_18 */

/* blackbox module Booth_Multiplier_bbox_17 */

/* blackbox module Booth_Multiplier_bbox_16 */

/* blackbox module Booth_Multiplier_bbox_15 */

/* blackbox module Booth_Multiplier_bbox_14 */

/* blackbox module Booth_Multiplier_bbox_13 */

/* blackbox module Booth_Multiplier_bbox_12 */

/* blackbox module Booth_Multiplier_bbox_11 */

/* blackbox module Booth_Multiplier_bbox_10 */

/* blackbox module Booth_Multiplier_bbox_9 */

/* blackbox module Booth_Multiplier_bbox_8 */

/* blackbox module Booth_Multiplier_bbox_7 */

/* blackbox module Booth_Multiplier_bbox_6 */

/* blackbox module Booth_Multiplier_bbox_5 */

/* blackbox module Booth_Multiplier_bbox_4 */

/* blackbox module Booth_Multiplier_bbox_3 */

/* blackbox module Booth_Multiplier_bbox_2 */

/* blackbox module Booth_Multiplier_bbox_1 */

/* blackbox module Booth_Multiplier_bbox_0 */

/* blackbox module Booth_Multiplier_bbox */

module conv(\window[0][0] , \window[0][1] , \window[0][2] , \window[0][3] , 
      \window[0][4] , \window[1][0] , \window[1][1] , \window[1][2] , 
      \window[1][3] , \window[1][4] , \window[2][0] , \window[2][1] , 
      \window[2][2] , \window[2][3] , \window[2][4] , \window[3][0] , 
      \window[3][1] , \window[3][2] , \window[3][3] , \window[3][4] , 
      \window[4][0] , \window[4][1] , \window[4][2] , \window[4][3] , 
      \window[4][4] , \filter[0][0] , \filter[0][1] , \filter[0][2] , 
      \filter[0][3] , \filter[0][4] , \filter[1][0] , \filter[1][1] , 
      \filter[1][2] , \filter[1][3] , \filter[1][4] , \filter[2][0] , 
      \filter[2][1] , \filter[2][2] , \filter[2][3] , \filter[2][4] , 
      \filter[3][0] , \filter[3][1] , \filter[3][2] , \filter[3][3] , 
      \filter[3][4] , \filter[4][0] , \filter[4][1] , \filter[4][2] , 
      \filter[4][3] , \filter[4][4] , start, convResult, finish);
   input [15:0]\window[0][0] ;
   input [15:0]\window[0][1] ;
   input [15:0]\window[0][2] ;
   input [15:0]\window[0][3] ;
   input [15:0]\window[0][4] ;
   input [15:0]\window[1][0] ;
   input [15:0]\window[1][1] ;
   input [15:0]\window[1][2] ;
   input [15:0]\window[1][3] ;
   input [15:0]\window[1][4] ;
   input [15:0]\window[2][0] ;
   input [15:0]\window[2][1] ;
   input [15:0]\window[2][2] ;
   input [15:0]\window[2][3] ;
   input [15:0]\window[2][4] ;
   input [15:0]\window[3][0] ;
   input [15:0]\window[3][1] ;
   input [15:0]\window[3][2] ;
   input [15:0]\window[3][3] ;
   input [15:0]\window[3][4] ;
   input [15:0]\window[4][0] ;
   input [15:0]\window[4][1] ;
   input [15:0]\window[4][2] ;
   input [15:0]\window[4][3] ;
   input [15:0]\window[4][4] ;
   input [15:0]\filter[0][0] ;
   input [15:0]\filter[0][1] ;
   input [15:0]\filter[0][2] ;
   input [15:0]\filter[0][3] ;
   input [15:0]\filter[0][4] ;
   input [15:0]\filter[1][0] ;
   input [15:0]\filter[1][1] ;
   input [15:0]\filter[1][2] ;
   input [15:0]\filter[1][3] ;
   input [15:0]\filter[1][4] ;
   input [15:0]\filter[2][0] ;
   input [15:0]\filter[2][1] ;
   input [15:0]\filter[2][2] ;
   input [15:0]\filter[2][3] ;
   input [15:0]\filter[2][4] ;
   input [15:0]\filter[3][0] ;
   input [15:0]\filter[3][1] ;
   input [15:0]\filter[3][2] ;
   input [15:0]\filter[3][3] ;
   input [15:0]\filter[3][4] ;
   input [15:0]\filter[4][0] ;
   input [15:0]\filter[4][1] ;
   input [15:0]\filter[4][2] ;
   input [15:0]\filter[4][3] ;
   input [15:0]\filter[4][4] ;
   input start;
   output [15:0]convResult;
   output finish;

   wire [31:0]\products[24] ;
   wire [31:0]\products[23] ;
   wire [31:0]\products[22] ;
   wire [31:0]\products[21] ;
   wire [31:0]\products[20] ;
   wire [31:0]\products[19] ;
   wire [31:0]\products[18] ;
   wire [31:0]\products[17] ;
   wire [31:0]\products[16] ;
   wire [31:0]\products[15] ;
   wire [31:0]\products[14] ;
   wire [31:0]\products[13] ;
   wire [31:0]\products[12] ;
   wire [31:0]\products[11] ;
   wire [31:0]\products[10] ;
   wire [31:0]\products[9] ;
   wire [31:0]\products[8] ;
   wire [31:0]\products[7] ;
   wire [31:0]\products[6] ;
   wire [31:0]\products[5] ;
   wire [31:0]\products[4] ;
   wire [31:0]\products[3] ;
   wire [31:0]\products[2] ;
   wire [31:0]\products[1] ;
   wire [31:0]\products[0] ;

   Booth_Multiplier_bbox_23 genblk1_4_genblk1_4_booth (.p_0(\window[4][4] ), 
      .p_1(\filter[4][4] ), .p_2(\products[24] ));
   Booth_Multiplier_bbox_22 genblk1_4_genblk1_3_booth (.p_0(\window[4][3] ), 
      .p_1(\filter[4][3] ), .p_2(\products[23] ));
   Booth_Multiplier_bbox_21 genblk1_4_genblk1_2_booth (.p_0(\window[4][2] ), 
      .p_1(\filter[4][2] ), .p_2(\products[22] ));
   Booth_Multiplier_bbox_20 genblk1_4_genblk1_1_booth (.p_0(\window[4][1] ), 
      .p_1(\filter[4][1] ), .p_2(\products[21] ));
   Booth_Multiplier_bbox_19 genblk1_4_genblk1_0_booth (.p_0(\window[4][0] ), 
      .p_1(\filter[4][0] ), .p_2(\products[20] ));
   Booth_Multiplier_bbox_18 genblk1_3_genblk1_4_booth (.p_0(\window[3][4] ), 
      .p_1(\filter[3][4] ), .p_2(\products[19] ));
   Booth_Multiplier_bbox_17 genblk1_3_genblk1_3_booth (.p_0(\window[3][3] ), 
      .p_1(\filter[3][3] ), .p_2(\products[18] ));
   Booth_Multiplier_bbox_16 genblk1_3_genblk1_2_booth (.p_0(\window[3][2] ), 
      .p_1(\filter[3][2] ), .p_2(\products[17] ));
   Booth_Multiplier_bbox_15 genblk1_3_genblk1_1_booth (.p_0(\window[3][1] ), 
      .p_1(\filter[3][1] ), .p_2(\products[16] ));
   Booth_Multiplier_bbox_14 genblk1_3_genblk1_0_booth (.p_0(\window[3][0] ), 
      .p_1(\filter[3][0] ), .p_2(\products[15] ));
   Booth_Multiplier_bbox_13 genblk1_2_genblk1_4_booth (.p_0(\window[2][4] ), 
      .p_1(\filter[2][4] ), .p_2(\products[14] ));
   Booth_Multiplier_bbox_12 genblk1_2_genblk1_3_booth (.p_0(\window[2][3] ), 
      .p_1(\filter[2][3] ), .p_2(\products[13] ));
   Booth_Multiplier_bbox_11 genblk1_2_genblk1_2_booth (.p_0(\window[2][2] ), 
      .p_1(\filter[2][2] ), .p_2(\products[12] ));
   Booth_Multiplier_bbox_10 genblk1_2_genblk1_1_booth (.p_0(\window[2][1] ), 
      .p_1(\filter[2][1] ), .p_2(\products[11] ));
   Booth_Multiplier_bbox_9 genblk1_2_genblk1_0_booth (.p_0(\window[2][0] ), 
      .p_1(\filter[2][0] ), .p_2(\products[10] ));
   Booth_Multiplier_bbox_8 genblk1_1_genblk1_4_booth (.p_0(\window[1][4] ), 
      .p_1(\filter[1][4] ), .p_2(\products[9] ));
   Booth_Multiplier_bbox_7 genblk1_1_genblk1_3_booth (.p_0(\window[1][3] ), 
      .p_1(\filter[1][3] ), .p_2(\products[8] ));
   Booth_Multiplier_bbox_6 genblk1_1_genblk1_2_booth (.p_0(\window[1][2] ), 
      .p_1(\filter[1][2] ), .p_2(\products[7] ));
   Booth_Multiplier_bbox_5 genblk1_1_genblk1_1_booth (.p_0(\window[1][1] ), 
      .p_1(\filter[1][1] ), .p_2(\products[6] ));
   Booth_Multiplier_bbox_4 genblk1_1_genblk1_0_booth (.p_0(\window[1][0] ), 
      .p_1(\filter[1][0] ), .p_2(\products[5] ));
   Booth_Multiplier_bbox_3 genblk1_0_genblk1_4_booth (.p_0(\window[0][4] ), 
      .p_1(\filter[0][4] ), .p_2(\products[4] ));
   Booth_Multiplier_bbox_2 genblk1_0_genblk1_3_booth (.p_0(\window[0][3] ), 
      .p_1(\filter[0][3] ), .p_2(\products[3] ));
   Booth_Multiplier_bbox_1 genblk1_0_genblk1_2_booth (.p_0(\window[0][2] ), 
      .p_1(\filter[0][2] ), .p_2(\products[2] ));
   Booth_Multiplier_bbox_0 genblk1_0_genblk1_1_booth (.p_0(\window[0][1] ), 
      .p_1(\filter[0][1] ), .p_2(\products[1] ));
   Booth_Multiplier_bbox genblk1_0_genblk1_0_booth (.p_0(\window[0][0] ), 
      .p_1(\filter[0][0] ), .p_2(\products[0] ));
endmodule

module datapath__0_1152(p_0, p_1);
   input [15:0]p_0;
   output [15:0]p_1;

   HA_X1 i_2 (.A(p_0[2]), .B(p_0[1]), .CO(n_1), .S(p_1[2]));
   HA_X1 i_3 (.A(p_0[3]), .B(n_1), .CO(n_2), .S(p_1[3]));
   HA_X1 i_4 (.A(p_0[4]), .B(n_2), .CO(n_3), .S(p_1[4]));
   HA_X1 i_5 (.A(p_0[5]), .B(n_3), .CO(n_4), .S(p_1[5]));
   HA_X1 i_6 (.A(p_0[6]), .B(n_4), .CO(n_5), .S(p_1[6]));
   HA_X1 i_7 (.A(p_0[7]), .B(n_5), .CO(n_6), .S(p_1[7]));
   HA_X1 i_8 (.A(p_0[8]), .B(n_6), .CO(n_7), .S(p_1[8]));
   HA_X1 i_9 (.A(p_0[9]), .B(n_7), .CO(n_8), .S(p_1[9]));
   HA_X1 i_10 (.A(p_0[10]), .B(n_8), .CO(n_9), .S(p_1[10]));
   HA_X1 i_11 (.A(p_0[11]), .B(n_9), .CO(n_10), .S(p_1[11]));
   HA_X1 i_12 (.A(p_0[12]), .B(n_10), .CO(n_11), .S(p_1[12]));
   HA_X1 i_13 (.A(p_0[13]), .B(n_11), .CO(n_12), .S(p_1[13]));
   HA_X1 i_14 (.A(p_0[14]), .B(n_12), .CO(n_0), .S(p_1[14]));
   XOR2_X1 i_0 (.A(p_0[15]), .B(n_0), .Z(p_1[15]));
   INV_X1 i_1 (.A(p_0[1]), .ZN(p_1[1]));
endmodule

module datapath__0_1158(featureMapSize, p_0, p_1);
   input [6:0]featureMapSize;
   input [15:0]p_0;
   output [15:0]p_1;

   HA_X1 i_0 (.A(featureMapSize[0]), .B(p_0[0]), .CO(n_0), .S(p_1[0]));
   FA_X1 i_1 (.A(featureMapSize[1]), .B(p_0[1]), .CI(n_0), .CO(n_1), .S(p_1[1]));
   FA_X1 i_2 (.A(featureMapSize[2]), .B(p_0[2]), .CI(n_1), .CO(n_2), .S(p_1[2]));
   FA_X1 i_3 (.A(featureMapSize[1]), .B(p_0[3]), .CI(n_2), .CO(n_3), .S(p_1[3]));
   HA_X1 i_4 (.A(p_0[4]), .B(n_3), .CO(n_4), .S(p_1[4]));
   FA_X1 i_5 (.A(featureMapSize[5]), .B(p_0[5]), .CI(n_4), .CO(n_5), .S(p_1[5]));
   HA_X1 i_6 (.A(p_0[6]), .B(n_5), .CO(n_6), .S(p_1[6]));
   HA_X1 i_7 (.A(p_0[7]), .B(n_6), .CO(n_7), .S(p_1[7]));
   HA_X1 i_8 (.A(p_0[8]), .B(n_7), .CO(n_8), .S(p_1[8]));
   HA_X1 i_9 (.A(p_0[9]), .B(n_8), .CO(n_9), .S(p_1[9]));
   HA_X1 i_10 (.A(p_0[10]), .B(n_9), .CO(n_10), .S(p_1[10]));
   HA_X1 i_11 (.A(p_0[11]), .B(n_10), .CO(n_11), .S(p_1[11]));
   HA_X1 i_12 (.A(p_0[12]), .B(n_11), .CO(n_12), .S(p_1[12]));
   HA_X1 i_13 (.A(p_0[13]), .B(n_12), .CO(n_13), .S(p_1[13]));
   HA_X1 i_14 (.A(p_0[14]), .B(n_13), .CO(n_14), .S(p_1[14]));
   XOR2_X1 i_15 (.A(p_0[15]), .B(n_14), .Z(p_1[15]));
endmodule

module datapath__0_1167(poolingWindowY, p_0);
   input [31:0]poolingWindowY;
   output [31:0]p_0;

   HA_X1 i_1 (.A(poolingWindowY[2]), .B(poolingWindowY[1]), .CO(n_0), .S(p_0[2]));
   HA_X1 i_2 (.A(poolingWindowY[3]), .B(n_0), .CO(n_1), .S(p_0[3]));
   HA_X1 i_3 (.A(poolingWindowY[4]), .B(n_1), .CO(n_2), .S(p_0[4]));
   HA_X1 i_4 (.A(poolingWindowY[5]), .B(n_2), .CO(n_3), .S(p_0[5]));
   HA_X1 i_5 (.A(poolingWindowY[6]), .B(n_3), .CO(n_4), .S(p_0[6]));
   HA_X1 i_6 (.A(poolingWindowY[7]), .B(n_4), .CO(n_5), .S(p_0[7]));
   HA_X1 i_7 (.A(poolingWindowY[8]), .B(n_5), .CO(n_6), .S(p_0[8]));
   HA_X1 i_8 (.A(poolingWindowY[9]), .B(n_6), .CO(n_7), .S(p_0[9]));
   HA_X1 i_9 (.A(poolingWindowY[10]), .B(n_7), .CO(n_8), .S(p_0[10]));
   HA_X1 i_10 (.A(poolingWindowY[11]), .B(n_8), .CO(n_9), .S(p_0[11]));
   HA_X1 i_11 (.A(poolingWindowY[12]), .B(n_9), .CO(n_10), .S(p_0[12]));
   HA_X1 i_12 (.A(poolingWindowY[13]), .B(n_10), .CO(n_11), .S(p_0[13]));
   HA_X1 i_13 (.A(poolingWindowY[14]), .B(n_11), .CO(n_12), .S(p_0[14]));
   HA_X1 i_14 (.A(poolingWindowY[15]), .B(n_12), .CO(n_13), .S(p_0[15]));
   HA_X1 i_15 (.A(poolingWindowY[16]), .B(n_13), .CO(n_14), .S(p_0[16]));
   HA_X1 i_16 (.A(poolingWindowY[17]), .B(n_14), .CO(n_15), .S(p_0[17]));
   HA_X1 i_17 (.A(poolingWindowY[18]), .B(n_15), .CO(n_16), .S(p_0[18]));
   HA_X1 i_18 (.A(poolingWindowY[19]), .B(n_16), .CO(n_17), .S(p_0[19]));
   HA_X1 i_19 (.A(poolingWindowY[20]), .B(n_17), .CO(n_18), .S(p_0[20]));
   HA_X1 i_20 (.A(poolingWindowY[21]), .B(n_18), .CO(n_19), .S(p_0[21]));
   HA_X1 i_21 (.A(poolingWindowY[22]), .B(n_19), .CO(n_20), .S(p_0[22]));
   HA_X1 i_22 (.A(poolingWindowY[23]), .B(n_20), .CO(n_21), .S(p_0[23]));
   HA_X1 i_23 (.A(poolingWindowY[24]), .B(n_21), .CO(n_22), .S(p_0[24]));
   HA_X1 i_24 (.A(poolingWindowY[25]), .B(n_22), .CO(n_23), .S(p_0[25]));
   HA_X1 i_25 (.A(poolingWindowY[26]), .B(n_23), .CO(n_24), .S(p_0[26]));
   HA_X1 i_26 (.A(poolingWindowY[27]), .B(n_24), .CO(n_25), .S(p_0[27]));
   HA_X1 i_27 (.A(poolingWindowY[28]), .B(n_25), .CO(n_26), .S(p_0[28]));
   HA_X1 i_28 (.A(poolingWindowY[29]), .B(n_26), .CO(n_27), .S(p_0[29]));
   HA_X1 i_29 (.A(poolingWindowY[30]), .B(n_27), .CO(n_28), .S(p_0[30]));
   XOR2_X1 i_0 (.A(poolingWindowY[31]), .B(n_28), .Z(p_0[31]));
   INV_X1 i_30 (.A(poolingWindowY[1]), .ZN(p_0[1]));
endmodule

module datapath__0_1172(poolingWindowX, p_0);
   input [31:0]poolingWindowX;
   output [31:0]p_0;

   HA_X1 i_1 (.A(poolingWindowX[2]), .B(poolingWindowX[1]), .CO(n_0), .S(p_0[2]));
   HA_X1 i_2 (.A(poolingWindowX[3]), .B(n_0), .CO(n_1), .S(p_0[3]));
   HA_X1 i_3 (.A(poolingWindowX[4]), .B(n_1), .CO(n_2), .S(p_0[4]));
   HA_X1 i_4 (.A(poolingWindowX[5]), .B(n_2), .CO(n_3), .S(p_0[5]));
   HA_X1 i_5 (.A(poolingWindowX[6]), .B(n_3), .CO(n_4), .S(p_0[6]));
   HA_X1 i_6 (.A(poolingWindowX[7]), .B(n_4), .CO(n_5), .S(p_0[7]));
   HA_X1 i_7 (.A(poolingWindowX[8]), .B(n_5), .CO(n_6), .S(p_0[8]));
   HA_X1 i_8 (.A(poolingWindowX[9]), .B(n_6), .CO(n_7), .S(p_0[9]));
   HA_X1 i_9 (.A(poolingWindowX[10]), .B(n_7), .CO(n_8), .S(p_0[10]));
   HA_X1 i_10 (.A(poolingWindowX[11]), .B(n_8), .CO(n_9), .S(p_0[11]));
   HA_X1 i_11 (.A(poolingWindowX[12]), .B(n_9), .CO(n_10), .S(p_0[12]));
   HA_X1 i_12 (.A(poolingWindowX[13]), .B(n_10), .CO(n_11), .S(p_0[13]));
   HA_X1 i_13 (.A(poolingWindowX[14]), .B(n_11), .CO(n_12), .S(p_0[14]));
   HA_X1 i_14 (.A(poolingWindowX[15]), .B(n_12), .CO(n_13), .S(p_0[15]));
   HA_X1 i_15 (.A(poolingWindowX[16]), .B(n_13), .CO(n_14), .S(p_0[16]));
   HA_X1 i_16 (.A(poolingWindowX[17]), .B(n_14), .CO(n_15), .S(p_0[17]));
   HA_X1 i_17 (.A(poolingWindowX[18]), .B(n_15), .CO(n_16), .S(p_0[18]));
   HA_X1 i_18 (.A(poolingWindowX[19]), .B(n_16), .CO(n_17), .S(p_0[19]));
   HA_X1 i_19 (.A(poolingWindowX[20]), .B(n_17), .CO(n_18), .S(p_0[20]));
   HA_X1 i_20 (.A(poolingWindowX[21]), .B(n_18), .CO(n_19), .S(p_0[21]));
   HA_X1 i_21 (.A(poolingWindowX[22]), .B(n_19), .CO(n_20), .S(p_0[22]));
   HA_X1 i_22 (.A(poolingWindowX[23]), .B(n_20), .CO(n_21), .S(p_0[23]));
   HA_X1 i_23 (.A(poolingWindowX[24]), .B(n_21), .CO(n_22), .S(p_0[24]));
   HA_X1 i_24 (.A(poolingWindowX[25]), .B(n_22), .CO(n_23), .S(p_0[25]));
   HA_X1 i_25 (.A(poolingWindowX[26]), .B(n_23), .CO(n_24), .S(p_0[26]));
   HA_X1 i_26 (.A(poolingWindowX[27]), .B(n_24), .CO(n_25), .S(p_0[27]));
   HA_X1 i_27 (.A(poolingWindowX[28]), .B(n_25), .CO(n_26), .S(p_0[28]));
   HA_X1 i_28 (.A(poolingWindowX[29]), .B(n_26), .CO(n_27), .S(p_0[29]));
   HA_X1 i_29 (.A(poolingWindowX[30]), .B(n_27), .CO(n_28), .S(p_0[30]));
   XOR2_X1 i_0 (.A(poolingWindowX[31]), .B(n_28), .Z(p_0[31]));
   INV_X1 i_30 (.A(poolingWindowX[1]), .ZN(p_0[1]));
endmodule

module datapath__0_1174(poolingCounter, p_0);
   input [31:0]poolingCounter;
   output [31:0]p_0;

   HA_X1 i_1 (.A(poolingCounter[1]), .B(poolingCounter[0]), .CO(n_0), .S(p_0[1]));
   HA_X1 i_2 (.A(poolingCounter[2]), .B(n_0), .CO(n_1), .S(p_0[2]));
   HA_X1 i_3 (.A(poolingCounter[3]), .B(n_1), .CO(n_2), .S(p_0[3]));
   HA_X1 i_4 (.A(poolingCounter[4]), .B(n_2), .CO(n_3), .S(p_0[4]));
   HA_X1 i_5 (.A(poolingCounter[5]), .B(n_3), .CO(n_4), .S(p_0[5]));
   HA_X1 i_6 (.A(poolingCounter[6]), .B(n_4), .CO(n_5), .S(p_0[6]));
   HA_X1 i_7 (.A(poolingCounter[7]), .B(n_5), .CO(n_6), .S(p_0[7]));
   HA_X1 i_8 (.A(poolingCounter[8]), .B(n_6), .CO(n_7), .S(p_0[8]));
   HA_X1 i_9 (.A(poolingCounter[9]), .B(n_7), .CO(n_8), .S(p_0[9]));
   HA_X1 i_10 (.A(poolingCounter[10]), .B(n_8), .CO(n_9), .S(p_0[10]));
   HA_X1 i_11 (.A(poolingCounter[11]), .B(n_9), .CO(n_10), .S(p_0[11]));
   HA_X1 i_12 (.A(poolingCounter[12]), .B(n_10), .CO(n_11), .S(p_0[12]));
   HA_X1 i_13 (.A(poolingCounter[13]), .B(n_11), .CO(n_12), .S(p_0[13]));
   HA_X1 i_14 (.A(poolingCounter[14]), .B(n_12), .CO(n_13), .S(p_0[14]));
   HA_X1 i_15 (.A(poolingCounter[15]), .B(n_13), .CO(n_14), .S(p_0[15]));
   HA_X1 i_16 (.A(poolingCounter[16]), .B(n_14), .CO(n_15), .S(p_0[16]));
   HA_X1 i_17 (.A(poolingCounter[17]), .B(n_15), .CO(n_16), .S(p_0[17]));
   HA_X1 i_18 (.A(poolingCounter[18]), .B(n_16), .CO(n_17), .S(p_0[18]));
   HA_X1 i_19 (.A(poolingCounter[19]), .B(n_17), .CO(n_18), .S(p_0[19]));
   HA_X1 i_20 (.A(poolingCounter[20]), .B(n_18), .CO(n_19), .S(p_0[20]));
   HA_X1 i_21 (.A(poolingCounter[21]), .B(n_19), .CO(n_20), .S(p_0[21]));
   HA_X1 i_22 (.A(poolingCounter[22]), .B(n_20), .CO(n_21), .S(p_0[22]));
   HA_X1 i_23 (.A(poolingCounter[23]), .B(n_21), .CO(n_22), .S(p_0[23]));
   HA_X1 i_24 (.A(poolingCounter[24]), .B(n_22), .CO(n_23), .S(p_0[24]));
   HA_X1 i_25 (.A(poolingCounter[25]), .B(n_23), .CO(n_24), .S(p_0[25]));
   HA_X1 i_26 (.A(poolingCounter[26]), .B(n_24), .CO(n_25), .S(p_0[26]));
   HA_X1 i_27 (.A(poolingCounter[27]), .B(n_25), .CO(n_26), .S(p_0[27]));
   HA_X1 i_28 (.A(poolingCounter[28]), .B(n_26), .CO(n_27), .S(p_0[28]));
   HA_X1 i_29 (.A(poolingCounter[29]), .B(n_27), .CO(n_28), .S(p_0[29]));
   HA_X1 i_30 (.A(poolingCounter[30]), .B(n_28), .CO(n_29), .S(p_0[30]));
   XOR2_X1 i_0 (.A(poolingCounter[31]), .B(n_29), .Z(p_0[31]));
endmodule

module CNN(start, reset, finish, clk);
   input start;
   input reset;
   output finish;
   input clk;

   wire Mem_finish;
   wire [15:0]\Mem_input_data[4][4] ;
   wire [15:0]\Mem_input_data[4][3] ;
   wire [15:0]\Mem_input_data[4][2] ;
   wire [15:0]\Mem_input_data[4][1] ;
   wire [15:0]\Mem_input_data[4][0] ;
   wire [15:0]\Mem_input_data[3][4] ;
   wire [15:0]\Mem_input_data[3][3] ;
   wire [15:0]\Mem_input_data[3][2] ;
   wire [15:0]\Mem_input_data[3][1] ;
   wire [15:0]\Mem_input_data[3][0] ;
   wire [15:0]\Mem_input_data[2][4] ;
   wire [15:0]\Mem_input_data[2][3] ;
   wire [15:0]\Mem_input_data[2][2] ;
   wire [15:0]\Mem_input_data[2][1] ;
   wire [15:0]\Mem_input_data[2][0] ;
   wire [15:0]\Mem_input_data[1][4] ;
   wire [15:0]\Mem_input_data[1][3] ;
   wire [15:0]\Mem_input_data[1][2] ;
   wire [15:0]\Mem_input_data[1][1] ;
   wire [15:0]\Mem_input_data[1][0] ;
   wire [15:0]\Mem_input_data[0][4] ;
   wire [15:0]\Mem_input_data[0][3] ;
   wire [15:0]\Mem_input_data[0][2] ;
   wire [15:0]\Mem_input_data[0][1] ;
   wire [15:0]\Mem_input_data[0][0] ;
   wire FB_bias_or_filter;
   wire [15:0]FB_index_filter;
   wire [15:0]\FB_filter[4][4] ;
   wire [15:0]\FB_filter[4][3] ;
   wire [15:0]\FB_filter[4][2] ;
   wire [15:0]\FB_filter[4][1] ;
   wire [15:0]\FB_filter[4][0] ;
   wire [15:0]\FB_filter[3][4] ;
   wire [15:0]\FB_filter[3][3] ;
   wire [15:0]\FB_filter[3][2] ;
   wire [15:0]\FB_filter[3][1] ;
   wire [15:0]\FB_filter[3][0] ;
   wire [15:0]\FB_filter[2][4] ;
   wire [15:0]\FB_filter[2][3] ;
   wire [15:0]\FB_filter[2][2] ;
   wire [15:0]\FB_filter[2][1] ;
   wire [15:0]\FB_filter[2][0] ;
   wire [15:0]\FB_filter[1][4] ;
   wire [15:0]\FB_filter[1][3] ;
   wire [15:0]\FB_filter[1][2] ;
   wire [15:0]\FB_filter[1][1] ;
   wire [15:0]\FB_filter[1][0] ;
   wire [15:0]\FB_filter[0][4] ;
   wire [15:0]\FB_filter[0][3] ;
   wire [15:0]\FB_filter[0][2] ;
   wire [15:0]\FB_filter[0][1] ;
   wire [15:0]\FB_filter[0][0] ;
   wire [15:0]\DMA_CNN_output_data[4][4] ;
   wire [15:0]\DMA_CNN_output_data[4][3] ;
   wire [15:0]\DMA_CNN_output_data[4][2] ;
   wire [15:0]\DMA_CNN_output_data[4][1] ;
   wire [15:0]\DMA_CNN_output_data[4][0] ;
   wire [15:0]\DMA_CNN_output_data[3][4] ;
   wire [15:0]\DMA_CNN_output_data[3][3] ;
   wire [15:0]\DMA_CNN_output_data[3][2] ;
   wire [15:0]\DMA_CNN_output_data[3][1] ;
   wire [15:0]\DMA_CNN_output_data[3][0] ;
   wire [15:0]\DMA_CNN_output_data[2][4] ;
   wire [15:0]\DMA_CNN_output_data[2][3] ;
   wire [15:0]\DMA_CNN_output_data[2][2] ;
   wire [15:0]\DMA_CNN_output_data[2][1] ;
   wire [15:0]\DMA_CNN_output_data[2][0] ;
   wire [15:0]\DMA_CNN_output_data[1][4] ;
   wire [15:0]\DMA_CNN_output_data[1][3] ;
   wire [15:0]\DMA_CNN_output_data[1][2] ;
   wire [15:0]\DMA_CNN_output_data[1][1] ;
   wire [15:0]\DMA_CNN_output_data[1][0] ;
   wire [15:0]\DMA_CNN_output_data[0][4] ;
   wire [15:0]\DMA_CNN_output_data[0][3] ;
   wire [15:0]\DMA_CNN_output_data[0][2] ;
   wire [15:0]\DMA_CNN_output_data[0][1] ;
   wire [15:0]\DMA_CNN_output_data[0][0] ;
   wire [15:0]\filter[4][4] ;
   wire [15:0]\filter[4][3] ;
   wire [15:0]\filter[4][2] ;
   wire [15:0]\filter[4][1] ;
   wire [15:0]\filter[4][0] ;
   wire [15:0]\filter[3][4] ;
   wire [15:0]\filter[3][3] ;
   wire [15:0]\filter[3][2] ;
   wire [15:0]\filter[3][1] ;
   wire [15:0]\filter[3][0] ;
   wire [15:0]\filter[2][4] ;
   wire [15:0]\filter[2][3] ;
   wire [15:0]\filter[2][2] ;
   wire [15:0]\filter[2][1] ;
   wire [15:0]\filter[2][0] ;
   wire [15:0]\filter[1][4] ;
   wire [15:0]\filter[1][3] ;
   wire [15:0]\filter[1][2] ;
   wire [15:0]\filter[1][1] ;
   wire [15:0]\filter[1][0] ;
   wire [15:0]\filter[0][4] ;
   wire [15:0]\filter[0][3] ;
   wire [15:0]\filter[0][2] ;
   wire [15:0]\filter[0][1] ;
   wire [15:0]\filter[0][0] ;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_219;
   wire n_0_220;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_230;
   wire n_0_231;
   wire n_0_232;
   wire n_0_233;
   wire n_0_234;
   wire n_0_235;
   wire n_0_236;
   wire n_0_237;
   wire n_0_238;
   wire n_0_239;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_248;
   wire n_0_249;
   wire n_0_284;
   wire n_0_285;
   wire n_0_286;
   wire n_0_287;
   wire n_0_288;
   wire n_0_289;
   wire n_0_290;
   wire n_0_291;
   wire n_0_292;
   wire n_0_293;
   wire n_0_294;
   wire n_0_295;
   wire n_0_296;
   wire n_0_297;
   wire n_0_298;
   wire n_0_299;
   wire n_0_300;
   wire n_0_301;
   wire n_0_302;
   wire n_0_303;
   wire n_0_304;
   wire n_0_305;
   wire n_0_306;
   wire n_0_307;
   wire n_0_308;
   wire n_0_309;
   wire n_0_310;
   wire n_0_311;
   wire n_0_312;
   wire n_0_313;
   wire n_0_314;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire DMA_start;
   wire [15:0]DMA_start_address;
   wire [31:0]poolingState;
   wire n_0_31;
   wire [31:0]layerCounter;
   wire poolingReset;
   wire [15:0]writeAdress;
   wire [15:0]readAdress;
   wire n_0_32;
   wire [31:0]poolingWindowY;
   wire n_0_33;
   wire [31:0]poolingCounter;
   wire n_0_34;
   wire [31:0]poolingWindowX;
   wire n_0_35;
   wire n_0_0_1;
   wire n_0_0_32;
   wire n_0_0_13;
   wire n_0_0_33;
   wire n_0_0_21;
   wire n_0_0_34;
   wire n_0_0_22;
   wire n_0_0_35;
   wire n_0_0_23;
   wire n_0_0_36;
   wire n_0_0_0;
   wire n_0_0_37;
   wire n_0_0_2;
   wire n_0_0_38;
   wire n_0_0_3;
   wire n_0_0_39;
   wire n_0_0_4;
   wire n_0_0_40;
   wire n_0_0_5;
   wire n_0_0_41;
   wire n_0_0_6;
   wire n_0_0_42;
   wire n_0_0_7;
   wire n_0_0_43;
   wire n_0_0_8;
   wire n_0_0_44;
   wire n_0_0_9;
   wire n_0_0_45;
   wire n_0_0_10;
   wire n_0_0_46;
   wire n_0_0_11;
   wire n_0_0_47;
   wire n_0_0_12;
   wire n_0_0_48;
   wire n_0_0_14;
   wire n_0_0_49;
   wire n_0_0_15;
   wire n_0_0_50;
   wire n_0_0_16;
   wire n_0_0_51;
   wire n_0_0_17;
   wire n_0_0_52;
   wire n_0_0_18;
   wire n_0_0_53;
   wire n_0_0_19;
   wire n_0_0_54;
   wire n_0_0_20;
   wire n_0_139;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_0_58;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_315;
   wire n_0_316;
   wire n_0_317;
   wire n_0_318;
   wire n_0_319;
   wire n_0_320;
   wire n_0_321;
   wire n_0_322;
   wire n_0_323;
   wire n_0_324;
   wire n_0_325;
   wire n_0_326;
   wire n_0_327;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_283;
   wire n_0_282;
   wire n_0_0_59;
   wire n_0_281;
   wire n_0_0_60;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_256;
   wire n_0_257;
   wire n_0_258;
   wire n_0_259;
   wire n_0_260;
   wire n_0_261;
   wire n_0_262;
   wire n_0_263;
   wire n_0_264;
   wire n_0_265;
   wire n_0_266;
   wire n_0_267;
   wire n_0_268;
   wire n_0_269;
   wire n_0_270;
   wire n_0_271;
   wire n_0_272;
   wire n_0_273;
   wire n_0_274;
   wire n_0_275;
   wire n_0_276;
   wire n_0_277;
   wire n_0_278;
   wire n_0_279;
   wire n_0_280;
   wire n_0_218;
   wire n_0_202;
   wire n_0_0_61;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_0_62;
   wire n_0_206;
   wire n_0_0_63;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_215;
   wire n_0_216;
   wire n_0_0_64;
   wire n_0_141;
   wire n_0_140;
   wire n_0_0_65;
   wire n_0_183;
   wire n_0_0_66;
   wire n_0_184;
   wire n_0_0_67;
   wire n_0_185;
   wire n_0_0_68;
   wire n_0_186;
   wire n_0_0_69;
   wire n_0_0_70;
   wire n_0_187;
   wire n_0_0_71;
   wire n_0_188;
   wire n_0_0_72;
   wire n_0_189;
   wire n_0_0_73;
   wire n_0_0_74;
   wire n_0_190;
   wire n_0_0_75;
   wire n_0_0_76;
   wire n_0_191;
   wire n_0_0_77;
   wire n_0_192;
   wire n_0_0_78;
   wire n_0_0_79;
   wire n_0_193;
   wire n_0_0_80;
   wire n_0_194;
   wire n_0_0_81;
   wire n_0_195;
   wire n_0_0_82;
   wire n_0_196;
   wire n_0_0_83;
   wire n_0_197;
   wire n_0_0_84;
   wire n_0_198;
   wire n_0_0_85;
   wire n_0_0_86;
   wire n_0_0_87;
   wire n_0_0_88;
   wire n_0_0_89;
   wire n_0_0_90;
   wire n_0_0_91;
   wire n_0_0_92;
   wire n_0_0_93;
   wire n_0_0_94;
   wire n_0_0_95;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_0_96;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_0_97;
   wire n_0_0_98;
   wire n_0_126;
   wire n_0_0_99;
   wire n_0_127;
   wire n_0_128;
   wire n_0_0_100;
   wire n_0_0_101;
   wire n_0_0_102;
   wire n_0_129;
   wire n_0_0_103;
   wire n_0_130;
   wire n_0_0_104;
   wire n_0_131;
   wire n_0_132;
   wire n_0_0_105;
   wire n_0_0_106;
   wire n_0_133;
   wire n_0_0_107;
   wire n_0_0_24;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_0_108;
   wire n_0_138;
   wire n_0_0_109;
   wire n_0_0_110;
   wire n_0_0_111;
   wire n_0_0_112;
   wire n_0_0_113;
   wire n_0_180;
   wire n_0_142;
   wire n_0_0_114;
   wire n_0_0_115;
   wire n_0_0_116;
   wire n_0_0_117;
   wire n_0_0_118;
   wire n_0_0_119;
   wire n_0_0_120;
   wire n_0_0_121;
   wire n_0_0_122;
   wire n_0_0_123;
   wire n_0_0_124;
   wire n_0_0_125;
   wire n_0_0_126;
   wire n_0_0_127;
   wire n_0_0_128;
   wire n_0_0_129;
   wire n_0_0_130;
   wire n_0_0_131;
   wire n_0_0_132;
   wire n_0_0_133;
   wire n_0_0_134;
   wire n_0_0_135;
   wire n_0_0_136;
   wire n_0_0_137;
   wire n_0_0_138;
   wire n_0_0_139;
   wire n_0_0_140;
   wire n_0_0_141;
   wire n_0_0_142;
   wire n_0_0_143;
   wire n_0_0_144;
   wire n_0_0_145;
   wire n_0_0_146;
   wire n_0_0_147;
   wire n_0_0_148;
   wire n_0_0_149;
   wire n_0_0_150;
   wire n_0_0_151;
   wire n_0_0_152;
   wire n_0_0_153;
   wire n_0_0_154;
   wire n_0_0_155;
   wire n_0_0_156;
   wire n_0_0_157;
   wire n_0_0_158;
   wire n_0_0_159;
   wire n_0_0_160;
   wire n_0_0_161;
   wire n_0_0_162;
   wire n_0_0_163;
   wire n_0_0_164;
   wire n_0_0_165;
   wire n_0_0_166;
   wire n_0_0_167;
   wire n_0_0_168;
   wire n_0_0_169;
   wire n_0_0_170;
   wire n_0_0_171;
   wire n_0_0_172;
   wire n_0_0_173;
   wire n_0_0_174;
   wire n_0_0_175;
   wire n_0_0_176;
   wire n_0_0_177;
   wire n_0_0_178;
   wire n_0_0_179;
   wire n_0_0_180;
   wire n_0_0_181;
   wire n_0_0_182;
   wire n_0_0_183;
   wire n_0_181;
   wire n_0_0_184;
   wire n_0_0_185;
   wire n_0_143;
   wire n_0_0_186;
   wire n_0_144;
   wire n_0_0_187;
   wire n_0_0_188;
   wire n_0_145;
   wire n_0_0_189;
   wire n_0_0_190;
   wire n_0_0_191;
   wire n_0_162;
   wire n_0_0_192;
   wire n_0_163;
   wire n_0_0_193;
   wire n_0_164;
   wire n_0_0_194;
   wire n_0_0_195;
   wire n_0_0_27;
   wire n_0_0_196;
   wire n_0_165;
   wire n_0_0_197;
   wire n_0_166;
   wire n_0_0_198;
   wire n_0_167;
   wire n_0_168;
   wire n_0_0_199;
   wire n_0_0_200;
   wire n_0_0_201;
   wire n_0_0_202;
   wire n_0_169;
   wire n_0_0_203;
   wire n_0_0_204;
   wire n_0_0_25;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_0_205;
   wire n_0_174;
   wire n_0_0_206;
   wire n_0_0_207;
   wire n_0_0_208;
   wire n_0_0_209;
   wire n_0_0_26;
   wire n_0_175;
   wire n_0_0_28;
   wire n_0_176;
   wire n_0_0_210;
   wire n_0_0_211;
   wire n_0_0_212;
   wire n_0_0_29;
   wire n_0_177;
   wire n_0_178;
   wire n_0_0_213;
   wire n_0_0_214;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_0_215;
   wire n_0_0_216;
   wire n_0_0_217;
   wire n_0_0_218;
   wire n_0_0_219;
   wire n_0_0_220;
   wire n_0_0_221;
   wire n_0_0_222;
   wire n_0_0_223;
   wire n_0_0_224;
   wire n_0_0_225;
   wire n_0_0_226;
   wire n_0_0_227;
   wire n_0_0_228;
   wire n_0_0_229;
   wire n_0_201;
   wire n_0_179;
   wire n_0_182;
   wire n_0_199;
   wire n_0_200;
   wire n_0_217;

   RAM RAM1 (.enable(), .clk(clk), .address(), .write(), .\output_data[0][0] (
      \Mem_input_data[0][0] ), .\output_data[0][1] (\Mem_input_data[0][1] ), 
      .\output_data[0][2] (\Mem_input_data[0][2] ), .\output_data[0][3] (
      \Mem_input_data[0][3] ), .\output_data[0][4] (\Mem_input_data[0][4] ), 
      .\output_data[1][0] (\Mem_input_data[1][0] ), .\output_data[1][1] (
      \Mem_input_data[1][1] ), .\output_data[1][2] (\Mem_input_data[1][2] ), 
      .\output_data[1][3] (\Mem_input_data[1][3] ), .\output_data[1][4] (
      \Mem_input_data[1][4] ), .\output_data[2][0] (\Mem_input_data[2][0] ), 
      .\output_data[2][1] (\Mem_input_data[2][1] ), .\output_data[2][2] (
      \Mem_input_data[2][2] ), .\output_data[2][3] (\Mem_input_data[2][3] ), 
      .\output_data[2][4] (\Mem_input_data[2][4] ), .\output_data[3][0] (
      \Mem_input_data[3][0] ), .\output_data[3][1] (\Mem_input_data[3][1] ), 
      .\output_data[3][2] (\Mem_input_data[3][2] ), .\output_data[3][3] (
      \Mem_input_data[3][3] ), .\output_data[3][4] (\Mem_input_data[3][4] ), 
      .\output_data[4][0] (\Mem_input_data[4][0] ), .\output_data[4][1] (
      \Mem_input_data[4][1] ), .\output_data[4][2] (\Mem_input_data[4][2] ), 
      .\output_data[4][3] (\Mem_input_data[4][3] ), .\output_data[4][4] (
      \Mem_input_data[4][4] ), .offset({uc_0, uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, 
      uc_7, uc_8, 1'b0, uc_9, 1'b0, uc_10, uc_11, uc_12, uc_13}), .input_data(), 
      .finish(Mem_finish));
   DMA DMA1 (.start(DMA_start), .reset(), .finish_read(), .clk(clk), .address(
      DMA_start_address), .offset(), .read_write_filter_bias({1'b0, 1'b0}), 
      .filter_number(), .\CNN_output_data[0][0] (\DMA_CNN_output_data[0][0] ), 
      .\CNN_output_data[0][1] (\DMA_CNN_output_data[0][1] ), 
      .\CNN_output_data[0][2] (\DMA_CNN_output_data[0][2] ), 
      .\CNN_output_data[0][3] (\DMA_CNN_output_data[0][3] ), 
      .\CNN_output_data[0][4] (\DMA_CNN_output_data[0][4] ), 
      .\CNN_output_data[1][0] (\DMA_CNN_output_data[1][0] ), 
      .\CNN_output_data[1][1] (\DMA_CNN_output_data[1][1] ), 
      .\CNN_output_data[1][2] (\DMA_CNN_output_data[1][2] ), 
      .\CNN_output_data[1][3] (\DMA_CNN_output_data[1][3] ), 
      .\CNN_output_data[1][4] (\DMA_CNN_output_data[1][4] ), 
      .\CNN_output_data[2][0] (\DMA_CNN_output_data[2][0] ), 
      .\CNN_output_data[2][1] (\DMA_CNN_output_data[2][1] ), 
      .\CNN_output_data[2][2] (\DMA_CNN_output_data[2][2] ), 
      .\CNN_output_data[2][3] (\DMA_CNN_output_data[2][3] ), 
      .\CNN_output_data[2][4] (\DMA_CNN_output_data[2][4] ), 
      .\CNN_output_data[3][0] (\DMA_CNN_output_data[3][0] ), 
      .\CNN_output_data[3][1] (\DMA_CNN_output_data[3][1] ), 
      .\CNN_output_data[3][2] (\DMA_CNN_output_data[3][2] ), 
      .\CNN_output_data[3][3] (\DMA_CNN_output_data[3][3] ), 
      .\CNN_output_data[3][4] (\DMA_CNN_output_data[3][4] ), 
      .\CNN_output_data[4][0] (\DMA_CNN_output_data[4][0] ), 
      .\CNN_output_data[4][1] (\DMA_CNN_output_data[4][1] ), 
      .\CNN_output_data[4][2] (\DMA_CNN_output_data[4][2] ), 
      .\CNN_output_data[4][3] (\DMA_CNN_output_data[4][3] ), 
      .\CNN_output_data[4][4] (\DMA_CNN_output_data[4][4] ), .CNN_input_data({
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0}), .RAM_address(), .RAM_offset(), .RAM_write(), 
      .RAM_output_data(), .\RAM_input_data[0][0] (\Mem_input_data[0][0] ), 
      .\RAM_input_data[0][1] (\Mem_input_data[0][1] ), .\RAM_input_data[0][2] (
      \Mem_input_data[0][2] ), .\RAM_input_data[0][3] (\Mem_input_data[0][3] ), 
      .\RAM_input_data[0][4] (\Mem_input_data[0][4] ), .\RAM_input_data[1][0] (
      \Mem_input_data[1][0] ), .\RAM_input_data[1][1] (\Mem_input_data[1][1] ), 
      .\RAM_input_data[1][2] (\Mem_input_data[1][2] ), .\RAM_input_data[1][3] (
      \Mem_input_data[1][3] ), .\RAM_input_data[1][4] (\Mem_input_data[1][4] ), 
      .\RAM_input_data[2][0] (\Mem_input_data[2][0] ), .\RAM_input_data[2][1] (
      \Mem_input_data[2][1] ), .\RAM_input_data[2][2] (\Mem_input_data[2][2] ), 
      .\RAM_input_data[2][3] (\Mem_input_data[2][3] ), .\RAM_input_data[2][4] (
      \Mem_input_data[2][4] ), .\RAM_input_data[3][0] (\Mem_input_data[3][0] ), 
      .\RAM_input_data[3][1] (\Mem_input_data[3][1] ), .\RAM_input_data[3][2] (
      \Mem_input_data[3][2] ), .\RAM_input_data[3][3] (\Mem_input_data[3][3] ), 
      .\RAM_input_data[3][4] (\Mem_input_data[3][4] ), .\RAM_input_data[4][0] (
      \Mem_input_data[4][0] ), .\RAM_input_data[4][1] (\Mem_input_data[4][1] ), 
      .\RAM_input_data[4][2] (\Mem_input_data[4][2] ), .\RAM_input_data[4][3] (
      \Mem_input_data[4][3] ), .\RAM_input_data[4][4] (\Mem_input_data[4][4] ), 
      .RAM_finish(Mem_finish), .RAM_enable(), .FB_write(), .\FB_filter[0][0] (
      \FB_filter[0][0] ), .\FB_filter[0][1] (\FB_filter[0][1] ), 
      .\FB_filter[0][2] (\FB_filter[0][2] ), .\FB_filter[0][3] (
      \FB_filter[0][3] ), .\FB_filter[0][4] (\FB_filter[0][4] ), 
      .\FB_filter[1][0] (\FB_filter[1][0] ), .\FB_filter[1][1] (
      \FB_filter[1][1] ), .\FB_filter[1][2] (\FB_filter[1][2] ), 
      .\FB_filter[1][3] (\FB_filter[1][3] ), .\FB_filter[1][4] (
      \FB_filter[1][4] ), .\FB_filter[2][0] (\FB_filter[2][0] ), 
      .\FB_filter[2][1] (\FB_filter[2][1] ), .\FB_filter[2][2] (
      \FB_filter[2][2] ), .\FB_filter[2][3] (\FB_filter[2][3] ), 
      .\FB_filter[2][4] (\FB_filter[2][4] ), .\FB_filter[3][0] (
      \FB_filter[3][0] ), .\FB_filter[3][1] (\FB_filter[3][1] ), 
      .\FB_filter[3][2] (\FB_filter[3][2] ), .\FB_filter[3][3] (
      \FB_filter[3][3] ), .\FB_filter[3][4] (\FB_filter[3][4] ), 
      .\FB_filter[4][0] (\FB_filter[4][0] ), .\FB_filter[4][1] (
      \FB_filter[4][1] ), .\FB_filter[4][2] (\FB_filter[4][2] ), 
      .\FB_filter[4][3] (\FB_filter[4][3] ), .\FB_filter[4][4] (
      \FB_filter[4][4] ), .FB_index_filter(FB_index_filter), .\FB_bias[0] (), 
      .\FB_bias[1] (), .\FB_bias[2] (), .\FB_bias[3] (), .\FB_bias[4] (), 
      .\FB_bias[5] (), .\FB_bias[6] (), .\FB_bias[7] (), .\FB_bias[8] (), 
      .\FB_bias[9] (), .\FB_bias[10] (), .\FB_bias[11] (), .\FB_bias[12] (), 
      .\FB_bias[13] (), .\FB_bias[14] (), .\FB_bias[15] (), .\FB_bias[16] (), 
      .\FB_bias[17] (), .\FB_bias[18] (), .\FB_bias[19] (), .\FB_bias[20] (), 
      .\FB_bias[21] (), .\FB_bias[22] (), .\FB_bias[23] (), .\FB_bias[24] (), 
      .\FB_bias[25] (), .\FB_bias[26] (), .\FB_bias[27] (), .\FB_bias[28] (), 
      .\FB_bias[29] (), .\FB_bias[30] (), .\FB_bias[31] (), .\FB_bias[32] (), 
      .\FB_bias[33] (), .\FB_bias[34] (), .\FB_bias[35] (), .\FB_bias[36] (), 
      .\FB_bias[37] (), .\FB_bias[38] (), .\FB_bias[39] (), .\FB_bias[40] (), 
      .\FB_bias[41] (), .\FB_bias[42] (), .\FB_bias[43] (), .\FB_bias[44] (), 
      .\FB_bias[45] (), .\FB_bias[46] (), .\FB_bias[47] (), .\FB_bias[48] (), 
      .\FB_bias[49] (), .\FB_bias[50] (), .\FB_bias[51] (), .\FB_bias[52] (), 
      .\FB_bias[53] (), .\FB_bias[54] (), .\FB_bias[55] (), .\FB_bias[56] (), 
      .\FB_bias[57] (), .\FB_bias[58] (), .\FB_bias[59] (), .\FB_bias[60] (), 
      .\FB_bias[61] (), .\FB_bias[62] (), .\FB_bias[63] (), .\FB_bias[64] (), 
      .\FB_bias[65] (), .\FB_bias[66] (), .\FB_bias[67] (), .\FB_bias[68] (), 
      .\FB_bias[69] (), .\FB_bias[70] (), .\FB_bias[71] (), .\FB_bias[72] (), 
      .\FB_bias[73] (), .\FB_bias[74] (), .\FB_bias[75] (), .\FB_bias[76] (), 
      .\FB_bias[77] (), .\FB_bias[78] (), .\FB_bias[79] (), .\FB_bias[80] (), 
      .\FB_bias[81] (), .\FB_bias[82] (), .\FB_bias[83] (), .\FB_bias[84] (), 
      .\FB_bias[85] (), .\FB_bias[86] (), .\FB_bias[87] (), .\FB_bias[88] (), 
      .\FB_bias[89] (), .\FB_bias[90] (), .\FB_bias[91] (), .\FB_bias[92] (), 
      .\FB_bias[93] (), .\FB_bias[94] (), .\FB_bias[95] (), .\FB_bias[96] (), 
      .\FB_bias[97] (), .\FB_bias[98] (), .\FB_bias[99] (), .\FB_bias[100] (), 
      .\FB_bias[101] (), .\FB_bias[102] (), .\FB_bias[103] (), .\FB_bias[104] (), 
      .\FB_bias[105] (), .\FB_bias[106] (), .\FB_bias[107] (), .\FB_bias[108] (), 
      .\FB_bias[109] (), .\FB_bias[110] (), .\FB_bias[111] (), .\FB_bias[112] (), 
      .\FB_bias[113] (), .\FB_bias[114] (), .\FB_bias[115] (), .\FB_bias[116] (), 
      .\FB_bias[117] (), .\FB_bias[118] (), .\FB_bias[119] (), 
      .FB_bias_or_filter(FB_bias_or_filter));
   Filter_Buffer_5x5 FILTER_BUFFER (.read(1'b0), .\input_filter[0][0] (
      \FB_filter[0][0] ), .\input_filter[0][1] (\FB_filter[0][1] ), 
      .\input_filter[0][2] (\FB_filter[0][2] ), .\input_filter[0][3] (
      \FB_filter[0][3] ), .\input_filter[0][4] (\FB_filter[0][4] ), 
      .\input_filter[1][0] (\FB_filter[1][0] ), .\input_filter[1][1] (
      \FB_filter[1][1] ), .\input_filter[1][2] (\FB_filter[1][2] ), 
      .\input_filter[1][3] (\FB_filter[1][3] ), .\input_filter[1][4] (
      \FB_filter[1][4] ), .\input_filter[2][0] (\FB_filter[2][0] ), 
      .\input_filter[2][1] (\FB_filter[2][1] ), .\input_filter[2][2] (
      \FB_filter[2][2] ), .\input_filter[2][3] (\FB_filter[2][3] ), 
      .\input_filter[2][4] (\FB_filter[2][4] ), .\input_filter[3][0] (
      \FB_filter[3][0] ), .\input_filter[3][1] (\FB_filter[3][1] ), 
      .\input_filter[3][2] (\FB_filter[3][2] ), .\input_filter[3][3] (
      \FB_filter[3][3] ), .\input_filter[3][4] (\FB_filter[3][4] ), 
      .\input_filter[4][0] (\FB_filter[4][0] ), .\input_filter[4][1] (
      \FB_filter[4][1] ), .\input_filter[4][2] (\FB_filter[4][2] ), 
      .\input_filter[4][3] (\FB_filter[4][3] ), .\input_filter[4][4] (
      \FB_filter[4][4] ), .finish(), .\output_filter[0][0] (\filter[0][0] ), 
      .\output_filter[0][1] (\filter[0][1] ), .\output_filter[0][2] (
      \filter[0][2] ), .\output_filter[0][3] (\filter[0][3] ), 
      .\output_filter[0][4] (\filter[0][4] ), .\output_filter[1][0] (
      \filter[1][0] ), .\output_filter[1][1] (\filter[1][1] ), 
      .\output_filter[1][2] (\filter[1][2] ), .\output_filter[1][3] (
      \filter[1][3] ), .\output_filter[1][4] (\filter[1][4] ), 
      .\output_filter[2][0] (\filter[2][0] ), .\output_filter[2][1] (
      \filter[2][1] ), .\output_filter[2][2] (\filter[2][2] ), 
      .\output_filter[2][3] (\filter[2][3] ), .\output_filter[2][4] (
      \filter[2][4] ), .\output_filter[3][0] (\filter[3][0] ), 
      .\output_filter[3][1] (\filter[3][1] ), .\output_filter[3][2] (
      \filter[3][2] ), .\output_filter[3][3] (\filter[3][3] ), 
      .\output_filter[3][4] (\filter[3][4] ), .\output_filter[4][0] (
      \filter[4][0] ), .\output_filter[4][1] (\filter[4][1] ), 
      .\output_filter[4][2] (\filter[4][2] ), .\output_filter[4][3] (
      \filter[4][3] ), .\output_filter[4][4] (\filter[4][4] ), .index_buffer(
      FB_index_filter), .index_bias({uc_14, uc_15, uc_16, uc_17, uc_18, uc_19, 
      uc_20, uc_21, uc_22, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), 
      .\input_bias[0] (), .\input_bias[1] (), .\input_bias[2] (), 
      .\input_bias[3] (), .\input_bias[4] (), .\input_bias[5] (), 
      .\input_bias[6] (), .\input_bias[7] (), .\input_bias[8] (), 
      .\input_bias[9] (), .\input_bias[10] (), .\input_bias[11] (), 
      .\input_bias[12] (), .\input_bias[13] (), .\input_bias[14] (), 
      .\input_bias[15] (), .\input_bias[16] (), .\input_bias[17] (), 
      .\input_bias[18] (), .\input_bias[19] (), .\input_bias[20] (), 
      .\input_bias[21] (), .\input_bias[22] (), .\input_bias[23] (), 
      .\input_bias[24] (), .\input_bias[25] (), .\input_bias[26] (), 
      .\input_bias[27] (), .\input_bias[28] (), .\input_bias[29] (), 
      .\input_bias[30] (), .\input_bias[31] (), .\input_bias[32] (), 
      .\input_bias[33] (), .\input_bias[34] (), .\input_bias[35] (), 
      .\input_bias[36] (), .\input_bias[37] (), .\input_bias[38] (), 
      .\input_bias[39] (), .\input_bias[40] (), .\input_bias[41] (), 
      .\input_bias[42] (), .\input_bias[43] (), .\input_bias[44] (), 
      .\input_bias[45] (), .\input_bias[46] (), .\input_bias[47] (), 
      .\input_bias[48] (), .\input_bias[49] (), .\input_bias[50] (), 
      .\input_bias[51] (), .\input_bias[52] (), .\input_bias[53] (), 
      .\input_bias[54] (), .\input_bias[55] (), .\input_bias[56] (), 
      .\input_bias[57] (), .\input_bias[58] (), .\input_bias[59] (), 
      .\input_bias[60] (), .\input_bias[61] (), .\input_bias[62] (), 
      .\input_bias[63] (), .\input_bias[64] (), .\input_bias[65] (), 
      .\input_bias[66] (), .\input_bias[67] (), .\input_bias[68] (), 
      .\input_bias[69] (), .\input_bias[70] (), .\input_bias[71] (), 
      .\input_bias[72] (), .\input_bias[73] (), .\input_bias[74] (), 
      .\input_bias[75] (), .\input_bias[76] (), .\input_bias[77] (), 
      .\input_bias[78] (), .\input_bias[79] (), .\input_bias[80] (), 
      .\input_bias[81] (), .\input_bias[82] (), .\input_bias[83] (), 
      .\input_bias[84] (), .\input_bias[85] (), .\input_bias[86] (), 
      .\input_bias[87] (), .\input_bias[88] (), .\input_bias[89] (), 
      .\input_bias[90] (), .\input_bias[91] (), .\input_bias[92] (), 
      .\input_bias[93] (), .\input_bias[94] (), .\input_bias[95] (), 
      .\input_bias[96] (), .\input_bias[97] (), .\input_bias[98] (), 
      .\input_bias[99] (), .\input_bias[100] (), .\input_bias[101] (), 
      .\input_bias[102] (), .\input_bias[103] (), .\input_bias[104] (), 
      .\input_bias[105] (), .\input_bias[106] (), .\input_bias[107] (), 
      .\input_bias[108] (), .\input_bias[109] (), .\input_bias[110] (), 
      .\input_bias[111] (), .\input_bias[112] (), .\input_bias[113] (), 
      .\input_bias[114] (), .\input_bias[115] (), .\input_bias[116] (), 
      .\input_bias[117] (), .\input_bias[118] (), .\input_bias[119] (), 
      .bias_or_filter(FB_bias_or_filter), .output_bias());
   conv CONV1 (.\window[0][0] (\DMA_CNN_output_data[0][0] ), .\window[0][1] (
      \DMA_CNN_output_data[0][1] ), .\window[0][2] (\DMA_CNN_output_data[0][2] ), 
      .\window[0][3] (\DMA_CNN_output_data[0][3] ), .\window[0][4] (
      \DMA_CNN_output_data[0][4] ), .\window[1][0] (\DMA_CNN_output_data[1][0] ), 
      .\window[1][1] (\DMA_CNN_output_data[1][1] ), .\window[1][2] (
      \DMA_CNN_output_data[1][2] ), .\window[1][3] (\DMA_CNN_output_data[1][3] ), 
      .\window[1][4] (\DMA_CNN_output_data[1][4] ), .\window[2][0] (
      \DMA_CNN_output_data[2][0] ), .\window[2][1] (\DMA_CNN_output_data[2][1] ), 
      .\window[2][2] (\DMA_CNN_output_data[2][2] ), .\window[2][3] (
      \DMA_CNN_output_data[2][3] ), .\window[2][4] (\DMA_CNN_output_data[2][4] ), 
      .\window[3][0] (\DMA_CNN_output_data[3][0] ), .\window[3][1] (
      \DMA_CNN_output_data[3][1] ), .\window[3][2] (\DMA_CNN_output_data[3][2] ), 
      .\window[3][3] (\DMA_CNN_output_data[3][3] ), .\window[3][4] (
      \DMA_CNN_output_data[3][4] ), .\window[4][0] (\DMA_CNN_output_data[4][0] ), 
      .\window[4][1] (\DMA_CNN_output_data[4][1] ), .\window[4][2] (
      \DMA_CNN_output_data[4][2] ), .\window[4][3] (\DMA_CNN_output_data[4][3] ), 
      .\window[4][4] (\DMA_CNN_output_data[4][4] ), .\filter[0][0] (
      \filter[0][0] ), .\filter[0][1] (\filter[0][1] ), .\filter[0][2] (
      \filter[0][2] ), .\filter[0][3] (\filter[0][3] ), .\filter[0][4] (
      \filter[0][4] ), .\filter[1][0] (\filter[1][0] ), .\filter[1][1] (
      \filter[1][1] ), .\filter[1][2] (\filter[1][2] ), .\filter[1][3] (
      \filter[1][3] ), .\filter[1][4] (\filter[1][4] ), .\filter[2][0] (
      \filter[2][0] ), .\filter[2][1] (\filter[2][1] ), .\filter[2][2] (
      \filter[2][2] ), .\filter[2][3] (\filter[2][3] ), .\filter[2][4] (
      \filter[2][4] ), .\filter[3][0] (\filter[3][0] ), .\filter[3][1] (
      \filter[3][1] ), .\filter[3][2] (\filter[3][2] ), .\filter[3][3] (
      \filter[3][3] ), .\filter[3][4] (\filter[3][4] ), .\filter[4][0] (
      \filter[4][0] ), .\filter[4][1] (\filter[4][1] ), .\filter[4][2] (
      \filter[4][2] ), .\filter[4][3] (\filter[4][3] ), .\filter[4][4] (
      \filter[4][4] ), .start(1'b0), .convResult(), .finish());
   DFF_X1 finishCNN_reg (.D(n_0_182), .CK(clk), .Q(finish), .QN());
   datapath__0_1152 i_0_22 (.p_0({n_0_138, n_0_137, n_0_136, n_0_135, n_0_134, 
      n_0_133, n_0_132, n_0_131, n_0_130, n_0_129, n_0_128, n_0_127, n_0_126, 
      n_0_125, n_0_124, uc_23}), .p_1({n_0_89, n_0_88, n_0_87, n_0_86, n_0_85, 
      n_0_84, n_0_83, n_0_82, n_0_81, n_0_80, n_0_79, n_0_78, n_0_77, n_0_76, 
      n_0_75, uc_24}));
   datapath__0_1158 i_0_28 (.featureMapSize({1'b0, n_0_178, 1'b0, uc_25, n_0_176, 
      n_0_177, n_0_175}), .p_0({n_0_174, n_0_173, n_0_172, n_0_171, n_0_170, 
      n_0_169, n_0_168, n_0_167, n_0_166, n_0_165, n_0_164, n_0_163, n_0_162, 
      n_0_145, n_0_144, n_0_143}), .p_1({n_0_161, n_0_160, n_0_159, n_0_158, 
      n_0_157, n_0_156, n_0_155, n_0_154, n_0_153, n_0_152, n_0_151, n_0_150, 
      n_0_149, n_0_148, n_0_147, n_0_146}));
   datapath__0_1167 i_0_37 (.poolingWindowY({poolingWindowY[31], 
      poolingWindowY[30], poolingWindowY[29], poolingWindowY[28], 
      poolingWindowY[27], poolingWindowY[26], poolingWindowY[25], 
      poolingWindowY[24], poolingWindowY[23], poolingWindowY[22], 
      poolingWindowY[21], poolingWindowY[20], poolingWindowY[19], 
      poolingWindowY[18], poolingWindowY[17], poolingWindowY[16], 
      poolingWindowY[15], poolingWindowY[14], poolingWindowY[13], 
      poolingWindowY[12], poolingWindowY[11], poolingWindowY[10], 
      poolingWindowY[9], poolingWindowY[8], poolingWindowY[7], poolingWindowY[6], 
      poolingWindowY[5], poolingWindowY[4], poolingWindowY[3], poolingWindowY[2], 
      poolingWindowY[1], uc_26}), .p_0({n_0_249, n_0_248, n_0_247, n_0_246, 
      n_0_245, n_0_244, n_0_243, n_0_242, n_0_241, n_0_240, n_0_239, n_0_238, 
      n_0_237, n_0_236, n_0_235, n_0_234, n_0_233, n_0_232, n_0_231, n_0_230, 
      n_0_229, n_0_228, n_0_227, n_0_226, n_0_225, n_0_224, n_0_223, n_0_222, 
      n_0_221, n_0_220, n_0_219, uc_27}));
   datapath__0_1172 i_0_42 (.poolingWindowX({poolingWindowX[31], 
      poolingWindowX[30], poolingWindowX[29], poolingWindowX[28], 
      poolingWindowX[27], poolingWindowX[26], poolingWindowX[25], 
      poolingWindowX[24], poolingWindowX[23], poolingWindowX[22], 
      poolingWindowX[21], poolingWindowX[20], poolingWindowX[19], 
      poolingWindowX[18], poolingWindowX[17], poolingWindowX[16], 
      poolingWindowX[15], poolingWindowX[14], poolingWindowX[13], 
      poolingWindowX[12], poolingWindowX[11], poolingWindowX[10], 
      poolingWindowX[9], poolingWindowX[8], poolingWindowX[7], poolingWindowX[6], 
      poolingWindowX[5], poolingWindowX[4], poolingWindowX[3], poolingWindowX[2], 
      poolingWindowX[1], uc_28}), .p_0({n_0_314, n_0_313, n_0_312, n_0_311, 
      n_0_310, n_0_309, n_0_308, n_0_307, n_0_306, n_0_305, n_0_304, n_0_303, 
      n_0_302, n_0_301, n_0_300, n_0_299, n_0_298, n_0_297, n_0_296, n_0_295, 
      n_0_294, n_0_293, n_0_292, n_0_291, n_0_290, n_0_289, n_0_288, n_0_287, 
      n_0_286, n_0_285, n_0_284, uc_29}));
   datapath__0_1174 i_0_44 (.poolingCounter(poolingCounter), .p_0({n_0_30, 
      n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, 
      n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, 
      n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2, 
      n_0_1, n_0_0, uc_30}));
   DFF_X1 DMA_start_reg (.D(n_0_199), .CK(clk), .Q(DMA_start), .QN());
   DFF_X1 \DMA_start_address_reg[15]  (.D(n_0_216), .CK(n_0_179), .Q(
      DMA_start_address[15]), .QN());
   DFF_X1 \DMA_start_address_reg[14]  (.D(n_0_215), .CK(n_0_179), .Q(
      DMA_start_address[14]), .QN());
   DFF_X1 \DMA_start_address_reg[13]  (.D(n_0_214), .CK(n_0_179), .Q(
      DMA_start_address[13]), .QN());
   DFF_X1 \DMA_start_address_reg[12]  (.D(n_0_213), .CK(n_0_179), .Q(
      DMA_start_address[12]), .QN());
   DFF_X1 \DMA_start_address_reg[11]  (.D(n_0_212), .CK(n_0_179), .Q(
      DMA_start_address[11]), .QN());
   DFF_X1 \DMA_start_address_reg[10]  (.D(n_0_211), .CK(n_0_179), .Q(
      DMA_start_address[10]), .QN());
   DFF_X1 \DMA_start_address_reg[9]  (.D(n_0_210), .CK(n_0_179), .Q(
      DMA_start_address[9]), .QN());
   DFF_X1 \DMA_start_address_reg[8]  (.D(n_0_209), .CK(n_0_179), .Q(
      DMA_start_address[8]), .QN());
   DFF_X1 \DMA_start_address_reg[7]  (.D(n_0_208), .CK(n_0_179), .Q(
      DMA_start_address[7]), .QN());
   DFF_X1 \DMA_start_address_reg[6]  (.D(n_0_207), .CK(n_0_179), .Q(
      DMA_start_address[6]), .QN());
   DFF_X1 \DMA_start_address_reg[5]  (.D(n_0_206), .CK(n_0_179), .Q(
      DMA_start_address[5]), .QN());
   DFF_X1 \DMA_start_address_reg[4]  (.D(n_0_205), .CK(n_0_179), .Q(
      DMA_start_address[4]), .QN());
   DFF_X1 \DMA_start_address_reg[3]  (.D(n_0_204), .CK(n_0_179), .Q(
      DMA_start_address[3]), .QN());
   DFF_X1 \DMA_start_address_reg[2]  (.D(n_0_203), .CK(n_0_179), .Q(
      DMA_start_address[2]), .QN());
   DFF_X1 \DMA_start_address_reg[1]  (.D(n_0_202), .CK(n_0_179), .Q(
      DMA_start_address[1]), .QN());
   DFF_X1 \DMA_start_address_reg[0]  (.D(n_0_201), .CK(n_0_179), .Q(
      DMA_start_address[0]), .QN());
   DFF_X1 \poolingState_reg[0]  (.D(n_0_200), .CK(clk), .Q(poolingState[0]), 
      .QN());
   CLKGATETST_X1 clk_gate_layerCounter_reg (.CK(clk), .E(n_0_281), .SE(1'b0), 
      .GCK(n_0_31));
   DFF_X1 \layerCounter_reg[31]  (.D(n_0_42), .CK(n_0_31), .Q(layerCounter[31]), 
      .QN());
   DFF_X1 \layerCounter_reg[2]  (.D(n_0_41), .CK(n_0_31), .Q(layerCounter[2]), 
      .QN());
   DFF_X1 \layerCounter_reg[1]  (.D(n_0_40), .CK(n_0_31), .Q(layerCounter[1]), 
      .QN());
   DFF_X1 \layerCounter_reg[0]  (.D(n_0_39), .CK(n_0_31), .Q(layerCounter[0]), 
      .QN());
   DFF_X1 poolingReset_reg (.D(n_0_217), .CK(clk), .Q(poolingReset), .QN());
   DFF_X1 \writeAdress_reg[15]  (.D(n_0_123), .CK(n_0_35), .Q(writeAdress[15]), 
      .QN());
   DFF_X1 \writeAdress_reg[14]  (.D(n_0_122), .CK(n_0_35), .Q(writeAdress[14]), 
      .QN());
   DFF_X1 \writeAdress_reg[13]  (.D(n_0_121), .CK(n_0_35), .Q(writeAdress[13]), 
      .QN());
   DFF_X1 \writeAdress_reg[12]  (.D(n_0_120), .CK(n_0_35), .Q(writeAdress[12]), 
      .QN());
   DFF_X1 \writeAdress_reg[11]  (.D(n_0_119), .CK(n_0_35), .Q(writeAdress[11]), 
      .QN());
   DFF_X1 \writeAdress_reg[10]  (.D(n_0_118), .CK(n_0_35), .Q(writeAdress[10]), 
      .QN());
   DFF_X1 \writeAdress_reg[9]  (.D(n_0_117), .CK(n_0_35), .Q(writeAdress[9]), 
      .QN());
   DFF_X1 \writeAdress_reg[8]  (.D(n_0_116), .CK(n_0_35), .Q(writeAdress[8]), 
      .QN());
   DFF_X1 \writeAdress_reg[7]  (.D(n_0_115), .CK(n_0_35), .Q(writeAdress[7]), 
      .QN());
   DFF_X1 \writeAdress_reg[6]  (.D(n_0_114), .CK(n_0_35), .Q(writeAdress[6]), 
      .QN());
   DFF_X1 \writeAdress_reg[5]  (.D(n_0_113), .CK(n_0_35), .Q(writeAdress[5]), 
      .QN());
   DFF_X1 \writeAdress_reg[4]  (.D(n_0_112), .CK(n_0_35), .Q(writeAdress[4]), 
      .QN());
   DFF_X1 \writeAdress_reg[3]  (.D(n_0_111), .CK(n_0_35), .Q(writeAdress[3]), 
      .QN());
   DFF_X1 \writeAdress_reg[2]  (.D(n_0_110), .CK(n_0_35), .Q(writeAdress[2]), 
      .QN());
   DFF_X1 \writeAdress_reg[1]  (.D(n_0_109), .CK(n_0_35), .Q(writeAdress[1]), 
      .QN());
   DFF_X1 \readAdress_reg[15]  (.D(n_0_198), .CK(n_0_35), .Q(readAdress[15]), 
      .QN());
   DFF_X1 \readAdress_reg[14]  (.D(n_0_197), .CK(n_0_35), .Q(readAdress[14]), 
      .QN());
   DFF_X1 \readAdress_reg[13]  (.D(n_0_196), .CK(n_0_35), .Q(readAdress[13]), 
      .QN());
   DFF_X1 \readAdress_reg[12]  (.D(n_0_195), .CK(n_0_35), .Q(readAdress[12]), 
      .QN());
   DFF_X1 \readAdress_reg[11]  (.D(n_0_194), .CK(n_0_35), .Q(readAdress[11]), 
      .QN());
   DFF_X1 \readAdress_reg[10]  (.D(n_0_193), .CK(n_0_35), .Q(readAdress[10]), 
      .QN());
   DFF_X1 \readAdress_reg[9]  (.D(n_0_192), .CK(n_0_35), .Q(readAdress[9]), 
      .QN());
   DFF_X1 \readAdress_reg[8]  (.D(n_0_191), .CK(n_0_35), .Q(readAdress[8]), 
      .QN());
   DFF_X1 \readAdress_reg[7]  (.D(n_0_190), .CK(n_0_35), .Q(readAdress[7]), 
      .QN());
   DFF_X1 \readAdress_reg[6]  (.D(n_0_189), .CK(n_0_35), .Q(readAdress[6]), 
      .QN());
   DFF_X1 \readAdress_reg[5]  (.D(n_0_188), .CK(n_0_35), .Q(readAdress[5]), 
      .QN());
   DFF_X1 \readAdress_reg[4]  (.D(n_0_187), .CK(n_0_35), .Q(readAdress[4]), 
      .QN());
   DFF_X1 \readAdress_reg[3]  (.D(n_0_186), .CK(n_0_35), .Q(readAdress[3]), 
      .QN());
   DFF_X1 \readAdress_reg[2]  (.D(n_0_185), .CK(n_0_35), .Q(readAdress[2]), 
      .QN());
   DFF_X1 \readAdress_reg[1]  (.D(n_0_184), .CK(n_0_35), .Q(readAdress[1]), 
      .QN());
   DFF_X1 \readAdress_reg[0]  (.D(n_0_183), .CK(n_0_35), .Q(readAdress[0]), 
      .QN());
   CLKGATETST_X1 clk_gate_poolingWindowY_reg (.CK(clk), .E(n_0_218), .SE(1'b0), 
      .GCK(n_0_32));
   DFF_X1 \poolingWindowY_reg[31]  (.D(n_0_280), .CK(n_0_32), .Q(
      poolingWindowY[31]), .QN());
   DFF_X1 \poolingWindowY_reg[30]  (.D(n_0_279), .CK(n_0_32), .Q(
      poolingWindowY[30]), .QN());
   DFF_X1 \poolingWindowY_reg[29]  (.D(n_0_278), .CK(n_0_32), .Q(
      poolingWindowY[29]), .QN());
   DFF_X1 \poolingWindowY_reg[28]  (.D(n_0_277), .CK(n_0_32), .Q(
      poolingWindowY[28]), .QN());
   DFF_X1 \poolingWindowY_reg[27]  (.D(n_0_276), .CK(n_0_32), .Q(
      poolingWindowY[27]), .QN());
   DFF_X1 \poolingWindowY_reg[26]  (.D(n_0_275), .CK(n_0_32), .Q(
      poolingWindowY[26]), .QN());
   DFF_X1 \poolingWindowY_reg[25]  (.D(n_0_274), .CK(n_0_32), .Q(
      poolingWindowY[25]), .QN());
   DFF_X1 \poolingWindowY_reg[24]  (.D(n_0_273), .CK(n_0_32), .Q(
      poolingWindowY[24]), .QN());
   DFF_X1 \poolingWindowY_reg[23]  (.D(n_0_272), .CK(n_0_32), .Q(
      poolingWindowY[23]), .QN());
   DFF_X1 \poolingWindowY_reg[22]  (.D(n_0_271), .CK(n_0_32), .Q(
      poolingWindowY[22]), .QN());
   DFF_X1 \poolingWindowY_reg[21]  (.D(n_0_270), .CK(n_0_32), .Q(
      poolingWindowY[21]), .QN());
   DFF_X1 \poolingWindowY_reg[20]  (.D(n_0_269), .CK(n_0_32), .Q(
      poolingWindowY[20]), .QN());
   DFF_X1 \poolingWindowY_reg[19]  (.D(n_0_268), .CK(n_0_32), .Q(
      poolingWindowY[19]), .QN());
   DFF_X1 \poolingWindowY_reg[18]  (.D(n_0_267), .CK(n_0_32), .Q(
      poolingWindowY[18]), .QN());
   DFF_X1 \poolingWindowY_reg[17]  (.D(n_0_266), .CK(n_0_32), .Q(
      poolingWindowY[17]), .QN());
   DFF_X1 \poolingWindowY_reg[16]  (.D(n_0_265), .CK(n_0_32), .Q(
      poolingWindowY[16]), .QN());
   DFF_X1 \poolingWindowY_reg[15]  (.D(n_0_264), .CK(n_0_32), .Q(
      poolingWindowY[15]), .QN());
   DFF_X1 \poolingWindowY_reg[14]  (.D(n_0_263), .CK(n_0_32), .Q(
      poolingWindowY[14]), .QN());
   DFF_X1 \poolingWindowY_reg[13]  (.D(n_0_262), .CK(n_0_32), .Q(
      poolingWindowY[13]), .QN());
   DFF_X1 \poolingWindowY_reg[12]  (.D(n_0_261), .CK(n_0_32), .Q(
      poolingWindowY[12]), .QN());
   DFF_X1 \poolingWindowY_reg[11]  (.D(n_0_260), .CK(n_0_32), .Q(
      poolingWindowY[11]), .QN());
   DFF_X1 \poolingWindowY_reg[10]  (.D(n_0_259), .CK(n_0_32), .Q(
      poolingWindowY[10]), .QN());
   DFF_X1 \poolingWindowY_reg[9]  (.D(n_0_258), .CK(n_0_32), .Q(
      poolingWindowY[9]), .QN());
   DFF_X1 \poolingWindowY_reg[8]  (.D(n_0_257), .CK(n_0_32), .Q(
      poolingWindowY[8]), .QN());
   DFF_X1 \poolingWindowY_reg[7]  (.D(n_0_256), .CK(n_0_32), .Q(
      poolingWindowY[7]), .QN());
   DFF_X1 \poolingWindowY_reg[6]  (.D(n_0_255), .CK(n_0_32), .Q(
      poolingWindowY[6]), .QN());
   DFF_X1 \poolingWindowY_reg[5]  (.D(n_0_254), .CK(n_0_32), .Q(
      poolingWindowY[5]), .QN());
   DFF_X1 \poolingWindowY_reg[4]  (.D(n_0_253), .CK(n_0_32), .Q(
      poolingWindowY[4]), .QN());
   DFF_X1 \poolingWindowY_reg[3]  (.D(n_0_252), .CK(n_0_32), .Q(
      poolingWindowY[3]), .QN());
   DFF_X1 \poolingWindowY_reg[2]  (.D(n_0_251), .CK(n_0_32), .Q(
      poolingWindowY[2]), .QN());
   DFF_X1 \poolingWindowY_reg[1]  (.D(n_0_250), .CK(n_0_32), .Q(
      poolingWindowY[1]), .QN());
   CLKGATETST_X1 clk_gate_poolingCounter_reg (.CK(clk), .E(n_0_282), .SE(1'b0), 
      .GCK(n_0_33));
   DFF_X1 \poolingCounter_reg[31]  (.D(n_0_74), .CK(n_0_33), .Q(
      poolingCounter[31]), .QN());
   DFF_X1 \poolingCounter_reg[30]  (.D(n_0_73), .CK(n_0_33), .Q(
      poolingCounter[30]), .QN());
   DFF_X1 \poolingCounter_reg[29]  (.D(n_0_72), .CK(n_0_33), .Q(
      poolingCounter[29]), .QN());
   DFF_X1 \poolingCounter_reg[28]  (.D(n_0_71), .CK(n_0_33), .Q(
      poolingCounter[28]), .QN());
   DFF_X1 \poolingCounter_reg[27]  (.D(n_0_70), .CK(n_0_33), .Q(
      poolingCounter[27]), .QN());
   DFF_X1 \poolingCounter_reg[26]  (.D(n_0_69), .CK(n_0_33), .Q(
      poolingCounter[26]), .QN());
   DFF_X1 \poolingCounter_reg[25]  (.D(n_0_68), .CK(n_0_33), .Q(
      poolingCounter[25]), .QN());
   DFF_X1 \poolingCounter_reg[24]  (.D(n_0_67), .CK(n_0_33), .Q(
      poolingCounter[24]), .QN());
   DFF_X1 \poolingCounter_reg[23]  (.D(n_0_66), .CK(n_0_33), .Q(
      poolingCounter[23]), .QN());
   DFF_X1 \poolingCounter_reg[22]  (.D(n_0_65), .CK(n_0_33), .Q(
      poolingCounter[22]), .QN());
   DFF_X1 \poolingCounter_reg[21]  (.D(n_0_64), .CK(n_0_33), .Q(
      poolingCounter[21]), .QN());
   DFF_X1 \poolingCounter_reg[20]  (.D(n_0_63), .CK(n_0_33), .Q(
      poolingCounter[20]), .QN());
   DFF_X1 \poolingCounter_reg[19]  (.D(n_0_62), .CK(n_0_33), .Q(
      poolingCounter[19]), .QN());
   DFF_X1 \poolingCounter_reg[18]  (.D(n_0_61), .CK(n_0_33), .Q(
      poolingCounter[18]), .QN());
   DFF_X1 \poolingCounter_reg[17]  (.D(n_0_60), .CK(n_0_33), .Q(
      poolingCounter[17]), .QN());
   DFF_X1 \poolingCounter_reg[16]  (.D(n_0_59), .CK(n_0_33), .Q(
      poolingCounter[16]), .QN());
   DFF_X1 \poolingCounter_reg[15]  (.D(n_0_58), .CK(n_0_33), .Q(
      poolingCounter[15]), .QN());
   DFF_X1 \poolingCounter_reg[14]  (.D(n_0_57), .CK(n_0_33), .Q(
      poolingCounter[14]), .QN());
   DFF_X1 \poolingCounter_reg[13]  (.D(n_0_56), .CK(n_0_33), .Q(
      poolingCounter[13]), .QN());
   DFF_X1 \poolingCounter_reg[12]  (.D(n_0_55), .CK(n_0_33), .Q(
      poolingCounter[12]), .QN());
   DFF_X1 \poolingCounter_reg[11]  (.D(n_0_54), .CK(n_0_33), .Q(
      poolingCounter[11]), .QN());
   DFF_X1 \poolingCounter_reg[10]  (.D(n_0_53), .CK(n_0_33), .Q(
      poolingCounter[10]), .QN());
   DFF_X1 \poolingCounter_reg[9]  (.D(n_0_52), .CK(n_0_33), .Q(poolingCounter[9]), 
      .QN());
   DFF_X1 \poolingCounter_reg[8]  (.D(n_0_51), .CK(n_0_33), .Q(poolingCounter[8]), 
      .QN());
   DFF_X1 \poolingCounter_reg[7]  (.D(n_0_50), .CK(n_0_33), .Q(poolingCounter[7]), 
      .QN());
   DFF_X1 \poolingCounter_reg[6]  (.D(n_0_49), .CK(n_0_33), .Q(poolingCounter[6]), 
      .QN());
   DFF_X1 \poolingCounter_reg[5]  (.D(n_0_48), .CK(n_0_33), .Q(poolingCounter[5]), 
      .QN());
   DFF_X1 \poolingCounter_reg[4]  (.D(n_0_47), .CK(n_0_33), .Q(poolingCounter[4]), 
      .QN());
   DFF_X1 \poolingCounter_reg[3]  (.D(n_0_46), .CK(n_0_33), .Q(poolingCounter[3]), 
      .QN());
   DFF_X1 \poolingCounter_reg[2]  (.D(n_0_45), .CK(n_0_33), .Q(poolingCounter[2]), 
      .QN());
   DFF_X1 \poolingCounter_reg[1]  (.D(n_0_44), .CK(n_0_33), .Q(poolingCounter[1]), 
      .QN());
   DFF_X1 \poolingCounter_reg[0]  (.D(n_0_43), .CK(n_0_33), .Q(poolingCounter[0]), 
      .QN());
   CLKGATETST_X1 clk_gate_poolingWindowX_reg (.CK(clk), .E(n_0_283), .SE(1'b0), 
      .GCK(n_0_34));
   DFF_X1 \poolingWindowX_reg[31]  (.D(n_0_107), .CK(n_0_34), .Q(
      poolingWindowX[31]), .QN());
   DFF_X1 \poolingWindowX_reg[30]  (.D(n_0_106), .CK(n_0_34), .Q(
      poolingWindowX[30]), .QN());
   DFF_X1 \poolingWindowX_reg[29]  (.D(n_0_105), .CK(n_0_34), .Q(
      poolingWindowX[29]), .QN());
   DFF_X1 \poolingWindowX_reg[28]  (.D(n_0_104), .CK(n_0_34), .Q(
      poolingWindowX[28]), .QN());
   DFF_X1 \poolingWindowX_reg[27]  (.D(n_0_103), .CK(n_0_34), .Q(
      poolingWindowX[27]), .QN());
   DFF_X1 \poolingWindowX_reg[26]  (.D(n_0_102), .CK(n_0_34), .Q(
      poolingWindowX[26]), .QN());
   DFF_X1 \poolingWindowX_reg[25]  (.D(n_0_101), .CK(n_0_34), .Q(
      poolingWindowX[25]), .QN());
   DFF_X1 \poolingWindowX_reg[24]  (.D(n_0_100), .CK(n_0_34), .Q(
      poolingWindowX[24]), .QN());
   DFF_X1 \poolingWindowX_reg[23]  (.D(n_0_99), .CK(n_0_34), .Q(
      poolingWindowX[23]), .QN());
   DFF_X1 \poolingWindowX_reg[22]  (.D(n_0_98), .CK(n_0_34), .Q(
      poolingWindowX[22]), .QN());
   DFF_X1 \poolingWindowX_reg[21]  (.D(n_0_97), .CK(n_0_34), .Q(
      poolingWindowX[21]), .QN());
   DFF_X1 \poolingWindowX_reg[20]  (.D(n_0_96), .CK(n_0_34), .Q(
      poolingWindowX[20]), .QN());
   DFF_X1 \poolingWindowX_reg[19]  (.D(n_0_95), .CK(n_0_34), .Q(
      poolingWindowX[19]), .QN());
   DFF_X1 \poolingWindowX_reg[18]  (.D(n_0_94), .CK(n_0_34), .Q(
      poolingWindowX[18]), .QN());
   DFF_X1 \poolingWindowX_reg[17]  (.D(n_0_93), .CK(n_0_34), .Q(
      poolingWindowX[17]), .QN());
   DFF_X1 \poolingWindowX_reg[16]  (.D(n_0_92), .CK(n_0_34), .Q(
      poolingWindowX[16]), .QN());
   DFF_X1 \poolingWindowX_reg[15]  (.D(n_0_91), .CK(n_0_34), .Q(
      poolingWindowX[15]), .QN());
   DFF_X1 \poolingWindowX_reg[14]  (.D(n_0_90), .CK(n_0_34), .Q(
      poolingWindowX[14]), .QN());
   DFF_X1 \poolingWindowX_reg[13]  (.D(n_0_327), .CK(n_0_34), .Q(
      poolingWindowX[13]), .QN());
   DFF_X1 \poolingWindowX_reg[12]  (.D(n_0_326), .CK(n_0_34), .Q(
      poolingWindowX[12]), .QN());
   DFF_X1 \poolingWindowX_reg[11]  (.D(n_0_325), .CK(n_0_34), .Q(
      poolingWindowX[11]), .QN());
   DFF_X1 \poolingWindowX_reg[10]  (.D(n_0_324), .CK(n_0_34), .Q(
      poolingWindowX[10]), .QN());
   DFF_X1 \poolingWindowX_reg[9]  (.D(n_0_323), .CK(n_0_34), .Q(
      poolingWindowX[9]), .QN());
   DFF_X1 \poolingWindowX_reg[8]  (.D(n_0_322), .CK(n_0_34), .Q(
      poolingWindowX[8]), .QN());
   DFF_X1 \poolingWindowX_reg[7]  (.D(n_0_321), .CK(n_0_34), .Q(
      poolingWindowX[7]), .QN());
   DFF_X1 \poolingWindowX_reg[6]  (.D(n_0_320), .CK(n_0_34), .Q(
      poolingWindowX[6]), .QN());
   DFF_X1 \poolingWindowX_reg[5]  (.D(n_0_319), .CK(n_0_34), .Q(
      poolingWindowX[5]), .QN());
   DFF_X1 \poolingWindowX_reg[4]  (.D(n_0_318), .CK(n_0_34), .Q(
      poolingWindowX[4]), .QN());
   DFF_X1 \poolingWindowX_reg[3]  (.D(n_0_317), .CK(n_0_34), .Q(
      poolingWindowX[3]), .QN());
   DFF_X1 \poolingWindowX_reg[2]  (.D(n_0_316), .CK(n_0_34), .Q(
      poolingWindowX[2]), .QN());
   DFF_X1 \poolingWindowX_reg[1]  (.D(n_0_315), .CK(n_0_34), .Q(
      poolingWindowX[1]), .QN());
   CLKGATETST_X1 clk_gate_writeAdress_reg (.CK(clk), .E(n_0_108), .SE(1'b0), 
      .GCK(n_0_35));
   HA_X1 i_0_0_0 (.A(layerCounter[2]), .B(n_0_0_30), .CO(n_0_0_1), .S());
   FA_X1 i_0_0_1 (.A(n_0_0_57), .B(n_0_0_26), .CI(n_0_0_28), .CO(n_0_0_13), 
      .S(n_0_0_32));
   FA_X1 i_0_0_2 (.A(n_0_0_28), .B(n_0_0_29), .CI(n_0_0_24), .CO(n_0_0_21), 
      .S(n_0_0_33));
   HA_X1 i_0_0_3 (.A(n_0_0_29), .B(n_0_0_21), .CO(n_0_0_22), .S(n_0_0_34));
   FA_X1 i_0_0_4 (.A(n_0_0_56), .B(n_0_0_29), .CI(n_0_0_22), .CO(n_0_0_23), 
      .S(n_0_0_35));
   FA_X1 i_0_0_5 (.A(n_0_0_55), .B(n_0_0_29), .CI(n_0_0_31), .CO(n_0_0_0), 
      .S(n_0_0_36));
   FA_X1 i_0_0_6 (.A(n_0_0_31), .B(n_0_0_27), .CI(n_0_0_25), .CO(n_0_0_2), 
      .S(n_0_0_37));
   HA_X1 i_0_0_7 (.A(n_0_0_27), .B(n_0_0_2), .CO(n_0_0_3), .S(n_0_0_38));
   FA_X1 i_0_0_8 (.A(n_0_0_137), .B(n_0_0_27), .CI(n_0_0_3), .CO(n_0_0_4), 
      .S(n_0_0_39));
   HA_X1 i_0_0_9 (.A(n_0_145), .B(n_0_144), .CO(n_0_0_5), .S(n_0_0_40));
   HA_X1 i_0_0_10 (.A(n_0_162), .B(n_0_0_5), .CO(n_0_0_6), .S(n_0_0_41));
   HA_X1 i_0_0_11 (.A(n_0_163), .B(n_0_0_6), .CO(n_0_0_7), .S(n_0_0_42));
   HA_X1 i_0_0_12 (.A(n_0_164), .B(n_0_0_7), .CO(n_0_0_8), .S(n_0_0_43));
   HA_X1 i_0_0_13 (.A(n_0_165), .B(n_0_0_8), .CO(n_0_0_9), .S(n_0_0_44));
   HA_X1 i_0_0_14 (.A(n_0_166), .B(n_0_0_9), .CO(n_0_0_10), .S(n_0_0_45));
   HA_X1 i_0_0_15 (.A(n_0_167), .B(n_0_0_10), .CO(n_0_0_11), .S(n_0_0_46));
   HA_X1 i_0_0_16 (.A(n_0_168), .B(n_0_0_11), .CO(n_0_0_12), .S(n_0_0_47));
   HA_X1 i_0_0_17 (.A(n_0_169), .B(n_0_0_12), .CO(n_0_0_14), .S(n_0_0_48));
   HA_X1 i_0_0_18 (.A(n_0_170), .B(n_0_0_14), .CO(n_0_0_15), .S(n_0_0_49));
   HA_X1 i_0_0_19 (.A(n_0_171), .B(n_0_0_15), .CO(n_0_0_16), .S(n_0_0_50));
   HA_X1 i_0_0_20 (.A(n_0_172), .B(n_0_0_16), .CO(n_0_0_17), .S(n_0_0_51));
   HA_X1 i_0_0_21 (.A(n_0_173), .B(n_0_0_17), .CO(n_0_0_18), .S(n_0_0_52));
   HA_X1 i_0_0_22 (.A(layerCounter[1]), .B(layerCounter[0]), .CO(n_0_0_19), 
      .S(n_0_0_53));
   HA_X1 i_0_0_23 (.A(layerCounter[2]), .B(n_0_0_19), .CO(n_0_0_20), .S(n_0_0_54));
   AND2_X1 i_0_0_24 (.A1(n_0_0_114), .A2(n_0_0_221), .ZN(n_0_139));
   NAND2_X1 i_0_0_25 (.A1(n_0_0_211), .A2(n_0_0_27), .ZN(n_0_0_55));
   NAND2_X1 i_0_0_26 (.A1(n_0_0_29), .A2(n_0_0_211), .ZN(n_0_0_56));
   OAI21_X1 i_0_0_27 (.A(n_0_0_29), .B1(n_0_0_101), .B2(layerCounter[2]), 
      .ZN(n_0_0_57));
   NOR2_X1 i_0_0_28 (.A1(n_0_0_185), .A2(reset), .ZN(n_0_36));
   NOR3_X1 i_0_0_29 (.A1(poolingState[0]), .A2(DMA_start), .A3(reset), .ZN(
      n_0_37));
   AOI21_X1 i_0_0_30 (.A(reset), .B1(n_0_0_222), .B2(n_0_0_223), .ZN(n_0_38));
   NOR2_X1 i_0_0_31 (.A1(layerCounter[0]), .A2(reset), .ZN(n_0_39));
   AND2_X1 i_0_0_32 (.A1(n_0_0_221), .A2(n_0_0_53), .ZN(n_0_40));
   AND2_X1 i_0_0_33 (.A1(n_0_0_221), .A2(n_0_0_54), .ZN(n_0_41));
   NOR2_X1 i_0_0_34 (.A1(n_0_0_58), .A2(reset), .ZN(n_0_42));
   XNOR2_X1 i_0_0_35 (.A(layerCounter[31]), .B(n_0_0_20), .ZN(n_0_0_58));
   NOR3_X1 i_0_0_36 (.A1(poolingCounter[0]), .A2(reset), .A3(n_0_0_119), 
      .ZN(n_0_43));
   AND2_X1 i_0_0_37 (.A1(n_0_0), .A2(n_0_140), .ZN(n_0_44));
   AND2_X1 i_0_0_38 (.A1(n_0_1), .A2(n_0_140), .ZN(n_0_45));
   AND2_X1 i_0_0_39 (.A1(n_0_2), .A2(n_0_140), .ZN(n_0_46));
   AND2_X1 i_0_0_40 (.A1(n_0_3), .A2(n_0_140), .ZN(n_0_47));
   AND2_X1 i_0_0_41 (.A1(n_0_4), .A2(n_0_140), .ZN(n_0_48));
   AND2_X1 i_0_0_42 (.A1(n_0_5), .A2(n_0_140), .ZN(n_0_49));
   AND2_X1 i_0_0_43 (.A1(n_0_6), .A2(n_0_140), .ZN(n_0_50));
   AND2_X1 i_0_0_44 (.A1(n_0_7), .A2(n_0_140), .ZN(n_0_51));
   AND2_X1 i_0_0_45 (.A1(n_0_8), .A2(n_0_140), .ZN(n_0_52));
   AND2_X1 i_0_0_46 (.A1(n_0_9), .A2(n_0_140), .ZN(n_0_53));
   AND2_X1 i_0_0_47 (.A1(n_0_10), .A2(n_0_140), .ZN(n_0_54));
   AND2_X1 i_0_0_48 (.A1(n_0_11), .A2(n_0_140), .ZN(n_0_55));
   AND2_X1 i_0_0_49 (.A1(n_0_12), .A2(n_0_140), .ZN(n_0_56));
   AND2_X1 i_0_0_50 (.A1(n_0_13), .A2(n_0_140), .ZN(n_0_57));
   AND2_X1 i_0_0_51 (.A1(n_0_14), .A2(n_0_140), .ZN(n_0_58));
   AND2_X1 i_0_0_52 (.A1(n_0_15), .A2(n_0_140), .ZN(n_0_59));
   AND2_X1 i_0_0_53 (.A1(n_0_16), .A2(n_0_140), .ZN(n_0_60));
   AND2_X1 i_0_0_54 (.A1(n_0_17), .A2(n_0_140), .ZN(n_0_61));
   AND2_X1 i_0_0_55 (.A1(n_0_18), .A2(n_0_140), .ZN(n_0_62));
   AND2_X1 i_0_0_56 (.A1(n_0_19), .A2(n_0_140), .ZN(n_0_63));
   AND2_X1 i_0_0_57 (.A1(n_0_20), .A2(n_0_140), .ZN(n_0_64));
   AND2_X1 i_0_0_58 (.A1(n_0_21), .A2(n_0_140), .ZN(n_0_65));
   AND2_X1 i_0_0_59 (.A1(n_0_22), .A2(n_0_140), .ZN(n_0_66));
   AND2_X1 i_0_0_60 (.A1(n_0_23), .A2(n_0_140), .ZN(n_0_67));
   AND2_X1 i_0_0_61 (.A1(n_0_24), .A2(n_0_140), .ZN(n_0_68));
   AND2_X1 i_0_0_62 (.A1(n_0_25), .A2(n_0_140), .ZN(n_0_69));
   AND2_X1 i_0_0_63 (.A1(n_0_26), .A2(n_0_140), .ZN(n_0_70));
   AND2_X1 i_0_0_64 (.A1(n_0_27), .A2(n_0_140), .ZN(n_0_71));
   AND2_X1 i_0_0_65 (.A1(n_0_28), .A2(n_0_140), .ZN(n_0_72));
   AND2_X1 i_0_0_66 (.A1(n_0_29), .A2(n_0_140), .ZN(n_0_73));
   AND2_X1 i_0_0_67 (.A1(n_0_30), .A2(n_0_140), .ZN(n_0_74));
   AND2_X1 i_0_0_68 (.A1(n_0_284), .A2(n_0_0_59), .ZN(n_0_315));
   AND2_X1 i_0_0_69 (.A1(n_0_285), .A2(n_0_0_59), .ZN(n_0_316));
   AND2_X1 i_0_0_70 (.A1(n_0_286), .A2(n_0_0_59), .ZN(n_0_317));
   AND2_X1 i_0_0_71 (.A1(n_0_287), .A2(n_0_0_59), .ZN(n_0_318));
   AND2_X1 i_0_0_72 (.A1(n_0_288), .A2(n_0_0_59), .ZN(n_0_319));
   AND2_X1 i_0_0_73 (.A1(n_0_289), .A2(n_0_0_59), .ZN(n_0_320));
   AND2_X1 i_0_0_74 (.A1(n_0_290), .A2(n_0_0_59), .ZN(n_0_321));
   AND2_X1 i_0_0_75 (.A1(n_0_291), .A2(n_0_0_59), .ZN(n_0_322));
   AND2_X1 i_0_0_76 (.A1(n_0_292), .A2(n_0_0_59), .ZN(n_0_323));
   AND2_X1 i_0_0_77 (.A1(n_0_293), .A2(n_0_0_59), .ZN(n_0_324));
   AND2_X1 i_0_0_78 (.A1(n_0_294), .A2(n_0_0_59), .ZN(n_0_325));
   AND2_X1 i_0_0_79 (.A1(n_0_295), .A2(n_0_0_59), .ZN(n_0_326));
   AND2_X1 i_0_0_80 (.A1(n_0_296), .A2(n_0_0_59), .ZN(n_0_327));
   AND2_X1 i_0_0_81 (.A1(n_0_297), .A2(n_0_0_59), .ZN(n_0_90));
   AND2_X1 i_0_0_82 (.A1(n_0_298), .A2(n_0_0_59), .ZN(n_0_91));
   AND2_X1 i_0_0_83 (.A1(n_0_299), .A2(n_0_0_59), .ZN(n_0_92));
   AND2_X1 i_0_0_84 (.A1(n_0_300), .A2(n_0_0_59), .ZN(n_0_93));
   AND2_X1 i_0_0_85 (.A1(n_0_301), .A2(n_0_0_59), .ZN(n_0_94));
   AND2_X1 i_0_0_86 (.A1(n_0_302), .A2(n_0_0_59), .ZN(n_0_95));
   AND2_X1 i_0_0_87 (.A1(n_0_303), .A2(n_0_0_59), .ZN(n_0_96));
   AND2_X1 i_0_0_88 (.A1(n_0_304), .A2(n_0_0_59), .ZN(n_0_97));
   AND2_X1 i_0_0_89 (.A1(n_0_305), .A2(n_0_0_59), .ZN(n_0_98));
   AND2_X1 i_0_0_90 (.A1(n_0_306), .A2(n_0_0_59), .ZN(n_0_99));
   AND2_X1 i_0_0_91 (.A1(n_0_307), .A2(n_0_0_59), .ZN(n_0_100));
   AND2_X1 i_0_0_92 (.A1(n_0_308), .A2(n_0_0_59), .ZN(n_0_101));
   AND2_X1 i_0_0_93 (.A1(n_0_309), .A2(n_0_0_59), .ZN(n_0_102));
   AND2_X1 i_0_0_94 (.A1(n_0_310), .A2(n_0_0_59), .ZN(n_0_103));
   AND2_X1 i_0_0_95 (.A1(n_0_311), .A2(n_0_0_59), .ZN(n_0_104));
   AND2_X1 i_0_0_96 (.A1(n_0_312), .A2(n_0_0_59), .ZN(n_0_105));
   AND2_X1 i_0_0_97 (.A1(n_0_313), .A2(n_0_0_59), .ZN(n_0_106));
   AND2_X1 i_0_0_98 (.A1(n_0_314), .A2(n_0_0_59), .ZN(n_0_107));
   AOI21_X1 i_0_0_99 (.A(n_0_0_113), .B1(n_0_0_115), .B2(n_0_0_221), .ZN(n_0_283));
   NOR2_X1 i_0_0_100 (.A1(n_0_0_65), .A2(n_0_0_59), .ZN(n_0_282));
   NOR3_X1 i_0_0_101 (.A1(reset), .A2(n_0_0_143), .A3(n_0_0_119), .ZN(n_0_0_59));
   INV_X1 i_0_0_102 (.A(n_0_0_60), .ZN(n_0_281));
   AOI21_X1 i_0_0_103 (.A(reset), .B1(n_0_0_117), .B2(n_0_0_183), .ZN(n_0_0_60));
   AND2_X1 i_0_0_104 (.A1(n_0_219), .A2(n_0_0_113), .ZN(n_0_250));
   AND2_X1 i_0_0_105 (.A1(n_0_220), .A2(n_0_0_113), .ZN(n_0_251));
   AND2_X1 i_0_0_106 (.A1(n_0_221), .A2(n_0_0_113), .ZN(n_0_252));
   AND2_X1 i_0_0_107 (.A1(n_0_222), .A2(n_0_0_113), .ZN(n_0_253));
   AND2_X1 i_0_0_108 (.A1(n_0_223), .A2(n_0_0_113), .ZN(n_0_254));
   AND2_X1 i_0_0_109 (.A1(n_0_224), .A2(n_0_0_113), .ZN(n_0_255));
   AND2_X1 i_0_0_110 (.A1(n_0_225), .A2(n_0_0_113), .ZN(n_0_256));
   AND2_X1 i_0_0_111 (.A1(n_0_226), .A2(n_0_0_113), .ZN(n_0_257));
   AND2_X1 i_0_0_112 (.A1(n_0_227), .A2(n_0_0_113), .ZN(n_0_258));
   AND2_X1 i_0_0_113 (.A1(n_0_228), .A2(n_0_0_113), .ZN(n_0_259));
   AND2_X1 i_0_0_114 (.A1(n_0_229), .A2(n_0_0_113), .ZN(n_0_260));
   AND2_X1 i_0_0_115 (.A1(n_0_230), .A2(n_0_0_113), .ZN(n_0_261));
   AND2_X1 i_0_0_116 (.A1(n_0_231), .A2(n_0_0_113), .ZN(n_0_262));
   AND2_X1 i_0_0_117 (.A1(n_0_232), .A2(n_0_0_113), .ZN(n_0_263));
   AND2_X1 i_0_0_118 (.A1(n_0_233), .A2(n_0_0_113), .ZN(n_0_264));
   AND2_X1 i_0_0_119 (.A1(n_0_234), .A2(n_0_0_113), .ZN(n_0_265));
   AND2_X1 i_0_0_120 (.A1(n_0_235), .A2(n_0_0_113), .ZN(n_0_266));
   AND2_X1 i_0_0_121 (.A1(n_0_236), .A2(n_0_0_113), .ZN(n_0_267));
   AND2_X1 i_0_0_122 (.A1(n_0_237), .A2(n_0_0_113), .ZN(n_0_268));
   AND2_X1 i_0_0_123 (.A1(n_0_238), .A2(n_0_0_113), .ZN(n_0_269));
   AND2_X1 i_0_0_124 (.A1(n_0_239), .A2(n_0_0_113), .ZN(n_0_270));
   AND2_X1 i_0_0_125 (.A1(n_0_240), .A2(n_0_0_113), .ZN(n_0_271));
   AND2_X1 i_0_0_126 (.A1(n_0_241), .A2(n_0_0_113), .ZN(n_0_272));
   AND2_X1 i_0_0_127 (.A1(n_0_242), .A2(n_0_0_113), .ZN(n_0_273));
   AND2_X1 i_0_0_128 (.A1(n_0_243), .A2(n_0_0_113), .ZN(n_0_274));
   AND2_X1 i_0_0_129 (.A1(n_0_244), .A2(n_0_0_113), .ZN(n_0_275));
   AND2_X1 i_0_0_130 (.A1(n_0_245), .A2(n_0_0_113), .ZN(n_0_276));
   AND2_X1 i_0_0_131 (.A1(n_0_246), .A2(n_0_0_113), .ZN(n_0_277));
   AND2_X1 i_0_0_132 (.A1(n_0_247), .A2(n_0_0_113), .ZN(n_0_278));
   AND2_X1 i_0_0_133 (.A1(n_0_248), .A2(n_0_0_113), .ZN(n_0_279));
   AND2_X1 i_0_0_134 (.A1(n_0_249), .A2(n_0_0_113), .ZN(n_0_280));
   OAI21_X1 i_0_0_135 (.A(n_0_0_221), .B1(n_0_0_116), .B2(n_0_0_94), .ZN(n_0_218));
   AOI21_X1 i_0_0_136 (.A(n_0_0_61), .B1(n_0_144), .B2(n_0_0_223), .ZN(n_0_202));
   NOR2_X1 i_0_0_137 (.A1(n_0_0_223), .A2(n_0_75), .ZN(n_0_0_61));
   MUX2_X1 i_0_0_138 (.A(n_0_0_40), .B(n_0_76), .S(poolingState[0]), .Z(n_0_203));
   MUX2_X1 i_0_0_139 (.A(n_0_0_41), .B(n_0_77), .S(poolingState[0]), .Z(n_0_204));
   OAI21_X1 i_0_0_140 (.A(n_0_0_62), .B1(n_0_0_216), .B2(poolingState[0]), 
      .ZN(n_0_205));
   NAND2_X1 i_0_0_141 (.A1(poolingState[0]), .A2(n_0_78), .ZN(n_0_0_62));
   OAI21_X1 i_0_0_142 (.A(n_0_0_63), .B1(n_0_0_215), .B2(poolingState[0]), 
      .ZN(n_0_206));
   NAND2_X1 i_0_0_143 (.A1(poolingState[0]), .A2(n_0_79), .ZN(n_0_0_63));
   MUX2_X1 i_0_0_144 (.A(n_0_0_44), .B(n_0_80), .S(poolingState[0]), .Z(n_0_207));
   MUX2_X1 i_0_0_145 (.A(n_0_0_45), .B(n_0_81), .S(poolingState[0]), .Z(n_0_208));
   MUX2_X1 i_0_0_146 (.A(n_0_0_46), .B(n_0_82), .S(poolingState[0]), .Z(n_0_209));
   MUX2_X1 i_0_0_147 (.A(n_0_0_47), .B(n_0_83), .S(poolingState[0]), .Z(n_0_210));
   MUX2_X1 i_0_0_148 (.A(n_0_0_48), .B(n_0_84), .S(poolingState[0]), .Z(n_0_211));
   MUX2_X1 i_0_0_149 (.A(n_0_0_49), .B(n_0_85), .S(poolingState[0]), .Z(n_0_212));
   MUX2_X1 i_0_0_150 (.A(n_0_0_50), .B(n_0_86), .S(poolingState[0]), .Z(n_0_213));
   MUX2_X1 i_0_0_151 (.A(n_0_0_51), .B(n_0_87), .S(poolingState[0]), .Z(n_0_214));
   MUX2_X1 i_0_0_152 (.A(n_0_0_52), .B(n_0_88), .S(poolingState[0]), .Z(n_0_215));
   AOI21_X1 i_0_0_153 (.A(n_0_0_64), .B1(n_0_0_90), .B2(n_0_0_223), .ZN(n_0_216));
   NOR2_X1 i_0_0_154 (.A1(n_0_0_223), .A2(n_0_89), .ZN(n_0_0_64));
   AOI21_X1 i_0_0_155 (.A(n_0_0_65), .B1(n_0_140), .B2(poolingReset), .ZN(
      n_0_141));
   NOR2_X1 i_0_0_156 (.A1(reset), .A2(n_0_0_119), .ZN(n_0_140));
   AOI21_X1 i_0_0_157 (.A(reset), .B1(n_0_0_183), .B2(layerCounter[0]), .ZN(
      n_0_0_65));
   AOI21_X1 i_0_0_158 (.A(n_0_0_66), .B1(n_0_0_94), .B2(n_0_0_186), .ZN(n_0_183));
   OAI21_X1 i_0_0_159 (.A(layerCounter[0]), .B1(n_0_0_94), .B2(n_0_146), 
      .ZN(n_0_0_66));
   OAI211_X1 i_0_0_160 (.A(n_0_0_67), .B(n_0_0_78), .C1(n_0_0_91), .C2(n_0_144), 
      .ZN(n_0_184));
   AOI22_X1 i_0_0_161 (.A1(n_0_147), .A2(n_0_0_93), .B1(n_0_0_87), .B2(
      readAdress[1]), .ZN(n_0_0_67));
   INV_X1 i_0_0_162 (.A(n_0_0_68), .ZN(n_0_185));
   AOI222_X1 i_0_0_163 (.A1(n_0_0_40), .A2(n_0_0_92), .B1(n_0_145), .B2(n_0_0_87), 
      .C1(n_0_148), .C2(n_0_0_93), .ZN(n_0_0_68));
   NAND3_X1 i_0_0_164 (.A1(n_0_0_69), .A2(n_0_0_70), .A3(n_0_0_78), .ZN(n_0_186));
   AOI22_X1 i_0_0_165 (.A1(n_0_149), .A2(n_0_0_93), .B1(n_0_0_87), .B2(
      readAdress[3]), .ZN(n_0_0_69));
   NAND2_X1 i_0_0_166 (.A1(n_0_0_41), .A2(n_0_0_92), .ZN(n_0_0_70));
   OAI21_X1 i_0_0_167 (.A(n_0_0_71), .B1(n_0_0_91), .B2(n_0_0_216), .ZN(n_0_187));
   AOI22_X1 i_0_0_168 (.A1(n_0_150), .A2(n_0_0_93), .B1(n_0_0_87), .B2(n_0_163), 
      .ZN(n_0_0_71));
   OAI21_X1 i_0_0_169 (.A(n_0_0_72), .B1(n_0_0_91), .B2(n_0_0_215), .ZN(n_0_188));
   AOI22_X1 i_0_0_170 (.A1(n_0_151), .A2(n_0_0_93), .B1(n_0_0_87), .B2(n_0_164), 
      .ZN(n_0_0_72));
   NAND3_X1 i_0_0_171 (.A1(n_0_0_73), .A2(n_0_0_74), .A3(n_0_0_78), .ZN(n_0_189));
   AOI22_X1 i_0_0_172 (.A1(n_0_152), .A2(n_0_0_93), .B1(n_0_0_87), .B2(
      readAdress[6]), .ZN(n_0_0_73));
   NAND2_X1 i_0_0_173 (.A1(n_0_0_44), .A2(n_0_0_92), .ZN(n_0_0_74));
   NAND3_X1 i_0_0_174 (.A1(n_0_0_75), .A2(n_0_0_76), .A3(n_0_0_78), .ZN(n_0_190));
   AOI22_X1 i_0_0_175 (.A1(n_0_0_45), .A2(n_0_0_92), .B1(n_0_0_87), .B2(
      readAdress[7]), .ZN(n_0_0_75));
   NAND2_X1 i_0_0_176 (.A1(n_0_153), .A2(n_0_0_93), .ZN(n_0_0_76));
   INV_X1 i_0_0_177 (.A(n_0_0_77), .ZN(n_0_191));
   AOI222_X1 i_0_0_178 (.A1(n_0_0_46), .A2(n_0_0_92), .B1(n_0_167), .B2(n_0_0_87), 
      .C1(n_0_154), .C2(n_0_0_93), .ZN(n_0_0_77));
   OAI21_X1 i_0_0_179 (.A(n_0_0_79), .B1(n_0_0_86), .B2(n_0_0_202), .ZN(n_0_192));
   OR2_X1 i_0_0_180 (.A1(n_0_0_86), .A2(poolingReset), .ZN(n_0_0_78));
   AOI22_X1 i_0_0_181 (.A1(n_0_155), .A2(n_0_0_93), .B1(n_0_0_92), .B2(n_0_0_47), 
      .ZN(n_0_0_79));
   OAI21_X1 i_0_0_182 (.A(n_0_0_80), .B1(n_0_0_86), .B2(n_0_0_203), .ZN(n_0_193));
   AOI22_X1 i_0_0_183 (.A1(n_0_156), .A2(n_0_0_93), .B1(n_0_0_92), .B2(n_0_0_48), 
      .ZN(n_0_0_80));
   INV_X1 i_0_0_184 (.A(n_0_0_81), .ZN(n_0_194));
   AOI222_X1 i_0_0_185 (.A1(n_0_0_49), .A2(n_0_0_92), .B1(n_0_170), .B2(n_0_0_87), 
      .C1(n_0_157), .C2(n_0_0_93), .ZN(n_0_0_81));
   INV_X1 i_0_0_186 (.A(n_0_0_82), .ZN(n_0_195));
   AOI222_X1 i_0_0_187 (.A1(n_0_0_50), .A2(n_0_0_92), .B1(n_0_171), .B2(n_0_0_87), 
      .C1(n_0_158), .C2(n_0_0_93), .ZN(n_0_0_82));
   INV_X1 i_0_0_188 (.A(n_0_0_83), .ZN(n_0_196));
   AOI222_X1 i_0_0_189 (.A1(n_0_0_51), .A2(n_0_0_92), .B1(n_0_172), .B2(n_0_0_87), 
      .C1(n_0_159), .C2(n_0_0_93), .ZN(n_0_0_83));
   OAI21_X1 i_0_0_190 (.A(n_0_0_84), .B1(n_0_0_86), .B2(n_0_0_205), .ZN(n_0_197));
   AOI22_X1 i_0_0_191 (.A1(n_0_160), .A2(n_0_0_93), .B1(n_0_0_92), .B2(n_0_0_52), 
      .ZN(n_0_0_84));
   OAI21_X1 i_0_0_192 (.A(n_0_0_85), .B1(n_0_0_90), .B2(n_0_0_91), .ZN(n_0_198));
   AOI22_X1 i_0_0_193 (.A1(n_0_161), .A2(n_0_0_93), .B1(n_0_0_87), .B2(n_0_174), 
      .ZN(n_0_0_85));
   NAND2_X1 i_0_0_194 (.A1(n_0_0_88), .A2(layerCounter[0]), .ZN(n_0_0_86));
   AOI21_X1 i_0_0_195 (.A(n_0_0_226), .B1(n_0_0_95), .B2(n_0_0_89), .ZN(n_0_0_87));
   NAND2_X1 i_0_0_196 (.A1(n_0_0_95), .A2(n_0_0_89), .ZN(n_0_0_88));
   OAI21_X1 i_0_0_197 (.A(n_0_0_164), .B1(DMA_start), .B2(poolingState[0]), 
      .ZN(n_0_0_89));
   XNOR2_X1 i_0_0_198 (.A(n_0_0_18), .B(n_0_174), .ZN(n_0_0_90));
   INV_X1 i_0_0_199 (.A(n_0_0_92), .ZN(n_0_0_91));
   NOR4_X1 i_0_0_200 (.A1(n_0_0_142), .A2(n_0_0_117), .A3(poolingState[0]), 
      .A4(DMA_start), .ZN(n_0_0_92));
   NOR2_X1 i_0_0_201 (.A1(n_0_0_226), .A2(n_0_0_94), .ZN(n_0_0_93));
   NAND2_X1 i_0_0_202 (.A1(n_0_0_163), .A2(n_0_0_95), .ZN(n_0_0_94));
   NOR2_X1 i_0_0_203 (.A1(n_0_0_143), .A2(n_0_0_119), .ZN(n_0_0_95));
   NOR2_X1 i_0_0_204 (.A1(n_0_0_116), .A2(reset), .ZN(n_0_108));
   AND2_X1 i_0_0_205 (.A1(layerCounter[0]), .A2(n_0_124), .ZN(n_0_109));
   AND2_X1 i_0_0_206 (.A1(n_0_125), .A2(layerCounter[0]), .ZN(n_0_110));
   AOI21_X1 i_0_0_207 (.A(n_0_0_96), .B1(poolingReset), .B2(n_0_0_218), .ZN(
      n_0_111));
   AOI21_X1 i_0_0_208 (.A(n_0_0_96), .B1(poolingReset), .B2(n_0_0_219), .ZN(
      n_0_112));
   AOI21_X1 i_0_0_209 (.A(n_0_0_96), .B1(poolingReset), .B2(n_0_0_220), .ZN(
      n_0_113));
   NAND2_X1 i_0_0_210 (.A1(n_0_0_190), .A2(layerCounter[0]), .ZN(n_0_0_96));
   OAI22_X1 i_0_0_211 (.A1(poolingReset), .A2(n_0_0_196), .B1(n_0_0_103), 
      .B2(n_0_0_226), .ZN(n_0_114));
   OAI22_X1 i_0_0_212 (.A1(poolingReset), .A2(n_0_0_196), .B1(n_0_0_104), 
      .B2(n_0_0_226), .ZN(n_0_115));
   AND2_X1 i_0_0_213 (.A1(n_0_131), .A2(layerCounter[0]), .ZN(n_0_116));
   AND2_X1 i_0_0_214 (.A1(n_0_132), .A2(layerCounter[0]), .ZN(n_0_117));
   AND2_X1 i_0_0_215 (.A1(n_0_133), .A2(layerCounter[0]), .ZN(n_0_118));
   AND2_X1 i_0_0_216 (.A1(n_0_134), .A2(layerCounter[0]), .ZN(n_0_119));
   AND2_X1 i_0_0_217 (.A1(n_0_135), .A2(layerCounter[0]), .ZN(n_0_120));
   AND2_X1 i_0_0_218 (.A1(n_0_136), .A2(layerCounter[0]), .ZN(n_0_121));
   AOI21_X1 i_0_0_219 (.A(n_0_0_226), .B1(n_0_0_110), .B2(n_0_0_108), .ZN(
      n_0_122));
   AOI21_X1 i_0_0_220 (.A(n_0_0_226), .B1(n_0_0_110), .B2(n_0_0_109), .ZN(
      n_0_123));
   AOI21_X1 i_0_0_221 (.A(n_0_0_191), .B1(poolingReset), .B2(n_0_0_217), 
      .ZN(n_0_124));
   OAI211_X1 i_0_0_222 (.A(n_0_0_98), .B(n_0_0_97), .C1(poolingReset), .C2(
      n_0_0_213), .ZN(n_0_125));
   NAND2_X1 i_0_0_223 (.A1(writeAdress[2]), .A2(poolingReset), .ZN(n_0_0_97));
   NAND2_X1 i_0_0_224 (.A1(n_0_0_102), .A2(n_0_0_200), .ZN(n_0_0_98));
   AOI21_X1 i_0_0_225 (.A(n_0_0_99), .B1(poolingReset), .B2(n_0_0_218), .ZN(
      n_0_126));
   NOR2_X1 i_0_0_226 (.A1(n_0_0_177), .A2(poolingReset), .ZN(n_0_0_99));
   AOI21_X1 i_0_0_227 (.A(n_0_0_100), .B1(poolingReset), .B2(n_0_0_219), 
      .ZN(n_0_127));
   AOI21_X1 i_0_0_228 (.A(n_0_0_100), .B1(poolingReset), .B2(n_0_0_220), 
      .ZN(n_0_128));
   NOR3_X1 i_0_0_229 (.A1(n_0_0_228), .A2(n_0_0_102), .A3(poolingReset), 
      .ZN(n_0_0_100));
   INV_X1 i_0_0_230 (.A(n_0_0_102), .ZN(n_0_0_101));
   NAND2_X1 i_0_0_231 (.A1(n_0_0_212), .A2(n_0_0_196), .ZN(n_0_0_102));
   OAI21_X1 i_0_0_232 (.A(n_0_0_103), .B1(n_0_0_28), .B2(poolingReset), .ZN(
      n_0_129));
   NAND2_X1 i_0_0_233 (.A1(writeAdress[6]), .A2(poolingReset), .ZN(n_0_0_103));
   OAI21_X1 i_0_0_234 (.A(n_0_0_104), .B1(n_0_0_28), .B2(poolingReset), .ZN(
      n_0_130));
   NAND2_X1 i_0_0_235 (.A1(writeAdress[7]), .A2(poolingReset), .ZN(n_0_0_104));
   MUX2_X1 i_0_0_236 (.A(n_0_0_32), .B(writeAdress[8]), .S(poolingReset), 
      .Z(n_0_131));
   OAI21_X1 i_0_0_237 (.A(n_0_0_106), .B1(n_0_0_105), .B2(poolingReset), 
      .ZN(n_0_132));
   XNOR2_X1 i_0_0_238 (.A(n_0_0_13), .B(n_0_0_177), .ZN(n_0_0_105));
   NAND2_X1 i_0_0_239 (.A1(writeAdress[9]), .A2(poolingReset), .ZN(n_0_0_106));
   OAI21_X1 i_0_0_240 (.A(n_0_0_107), .B1(n_0_0_24), .B2(poolingReset), .ZN(
      n_0_133));
   NAND2_X1 i_0_0_241 (.A1(writeAdress[10]), .A2(poolingReset), .ZN(n_0_0_107));
   AND2_X1 i_0_0_242 (.A1(n_0_0_177), .A2(n_0_0_13), .ZN(n_0_0_24));
   MUX2_X1 i_0_0_243 (.A(n_0_0_33), .B(writeAdress[11]), .S(poolingReset), 
      .Z(n_0_134));
   MUX2_X1 i_0_0_244 (.A(n_0_0_34), .B(writeAdress[12]), .S(poolingReset), 
      .Z(n_0_135));
   MUX2_X1 i_0_0_245 (.A(n_0_0_35), .B(writeAdress[13]), .S(poolingReset), 
      .Z(n_0_136));
   NAND2_X1 i_0_0_246 (.A1(n_0_0_110), .A2(n_0_0_108), .ZN(n_0_137));
   NAND2_X1 i_0_0_247 (.A1(writeAdress[14]), .A2(poolingReset), .ZN(n_0_0_108));
   NAND2_X1 i_0_0_248 (.A1(n_0_0_110), .A2(n_0_0_109), .ZN(n_0_138));
   NAND2_X1 i_0_0_249 (.A1(writeAdress[15]), .A2(poolingReset), .ZN(n_0_0_109));
   OAI21_X1 i_0_0_250 (.A(n_0_0_111), .B1(n_0_0_112), .B2(n_0_0_23), .ZN(
      n_0_0_110));
   AOI21_X1 i_0_0_251 (.A(poolingReset), .B1(n_0_0_23), .B2(n_0_0_112), .ZN(
      n_0_0_111));
   OAI21_X1 i_0_0_252 (.A(layerCounter[1]), .B1(n_0_0_228), .B2(layerCounter[0]), 
      .ZN(n_0_0_112));
   NOR2_X1 i_0_0_253 (.A1(n_0_0_142), .A2(reset), .ZN(n_0_0_113));
   OR2_X1 i_0_0_254 (.A1(reset), .A2(n_0_0_114), .ZN(n_0_180));
   OAI21_X1 i_0_0_255 (.A(n_0_0_221), .B1(n_0_0_142), .B2(n_0_0_115), .ZN(
      n_0_142));
   NOR3_X1 i_0_0_256 (.A1(n_0_0_115), .A2(poolingState[0]), .A3(n_0_0_142), 
      .ZN(n_0_0_114));
   NAND3_X1 i_0_0_257 (.A1(n_0_0_118), .A2(n_0_0_183), .A3(layerCounter[0]), 
      .ZN(n_0_0_115));
   NAND2_X1 i_0_0_258 (.A1(layerCounter[0]), .A2(n_0_0_183), .ZN(n_0_0_116));
   NAND2_X1 i_0_0_259 (.A1(n_0_0_118), .A2(layerCounter[0]), .ZN(n_0_0_117));
   INV_X1 i_0_0_260 (.A(n_0_0_119), .ZN(n_0_0_118));
   AOI21_X1 i_0_0_261 (.A(poolingCounter[31]), .B1(n_0_0_132), .B2(n_0_0_120), 
      .ZN(n_0_0_119));
   AND2_X1 i_0_0_262 (.A1(n_0_0_125), .A2(n_0_0_121), .ZN(n_0_0_120));
   NOR4_X1 i_0_0_263 (.A1(n_0_0_122), .A2(poolingCounter[28]), .A3(n_0_0_128), 
      .A4(poolingCounter[27]), .ZN(n_0_0_121));
   NAND4_X1 i_0_0_264 (.A1(n_0_0_126), .A2(n_0_0_124), .A3(n_0_0_123), .A4(
      n_0_0_127), .ZN(n_0_0_122));
   NOR4_X1 i_0_0_265 (.A1(poolingCounter[24]), .A2(poolingCounter[23]), .A3(
      poolingCounter[21]), .A4(poolingCounter[18]), .ZN(n_0_0_123));
   NOR2_X1 i_0_0_266 (.A1(poolingCounter[29]), .A2(poolingCounter[26]), .ZN(
      n_0_0_124));
   NOR4_X1 i_0_0_267 (.A1(poolingCounter[25]), .A2(poolingCounter[22]), .A3(
      poolingCounter[20]), .A4(poolingCounter[19]), .ZN(n_0_0_125));
   NOR2_X1 i_0_0_268 (.A1(poolingCounter[31]), .A2(poolingCounter[30]), .ZN(
      n_0_0_126));
   OAI21_X1 i_0_0_269 (.A(n_0_0_27), .B1(poolingCounter[5]), .B2(
      poolingCounter[6]), .ZN(n_0_0_127));
   NAND3_X1 i_0_0_270 (.A1(n_0_0_131), .A2(n_0_0_130), .A3(n_0_0_129), .ZN(
      n_0_0_128));
   NOR4_X1 i_0_0_271 (.A1(poolingCounter[17]), .A2(poolingCounter[14]), .A3(
      poolingCounter[12]), .A4(poolingCounter[11]), .ZN(n_0_0_129));
   NOR4_X1 i_0_0_272 (.A1(poolingCounter[16]), .A2(poolingCounter[15]), .A3(
      poolingCounter[13]), .A4(poolingCounter[10]), .ZN(n_0_0_130));
   NOR3_X1 i_0_0_273 (.A1(poolingCounter[9]), .A2(poolingCounter[8]), .A3(
      poolingCounter[7]), .ZN(n_0_0_131));
   OAI221_X1 i_0_0_274 (.A(n_0_0_134), .B1(n_0_0_133), .B2(n_0_0_27), .C1(
      n_0_0_136), .C2(poolingCounter[4]), .ZN(n_0_0_132));
   AND2_X1 i_0_0_275 (.A1(poolingCounter[6]), .A2(poolingCounter[5]), .ZN(
      n_0_0_133));
   OAI21_X1 i_0_0_276 (.A(n_0_0_135), .B1(n_0_0_140), .B2(n_0_0_138), .ZN(
      n_0_0_134));
   AOI21_X1 i_0_0_277 (.A(poolingCounter[3]), .B1(n_0_0_136), .B2(
      poolingCounter[4]), .ZN(n_0_0_135));
   INV_X1 i_0_0_278 (.A(n_0_0_137), .ZN(n_0_0_136));
   OAI21_X1 i_0_0_279 (.A(n_0_0_26), .B1(layerCounter[1]), .B2(n_0_0_228), 
      .ZN(n_0_0_137));
   OAI21_X1 i_0_0_280 (.A(n_0_0_27), .B1(n_0_0_210), .B2(n_0_0_139), .ZN(
      n_0_0_138));
   AND2_X1 i_0_0_281 (.A1(poolingCounter[2]), .A2(poolingCounter[1]), .ZN(
      n_0_0_139));
   AOI211_X1 i_0_0_282 (.A(poolingCounter[2]), .B(poolingCounter[1]), .C1(
      n_0_0_196), .C2(n_0_0_141), .ZN(n_0_0_140));
   NAND2_X1 i_0_0_283 (.A1(n_0_0_214), .A2(n_0_0_224), .ZN(n_0_0_141));
   OR2_X1 i_0_0_284 (.A1(n_0_0_163), .A2(n_0_0_143), .ZN(n_0_0_142));
   AOI21_X1 i_0_0_285 (.A(poolingWindowX[31]), .B1(n_0_0_144), .B2(n_0_0_158), 
      .ZN(n_0_0_143));
   INV_X1 i_0_0_286 (.A(n_0_0_145), .ZN(n_0_0_144));
   OR3_X1 i_0_0_287 (.A1(n_0_0_154), .A2(n_0_0_151), .A3(n_0_0_146), .ZN(
      n_0_0_145));
   NAND3_X1 i_0_0_288 (.A1(n_0_0_150), .A2(n_0_0_149), .A3(n_0_0_147), .ZN(
      n_0_0_146));
   AND2_X1 i_0_0_289 (.A1(n_0_0_148), .A2(n_0_0_177), .ZN(n_0_0_147));
   NOR4_X1 i_0_0_290 (.A1(poolingWindowX[8]), .A2(poolingWindowX[7]), .A3(
      poolingWindowX[6]), .A4(poolingWindowX[5]), .ZN(n_0_0_148));
   NOR4_X1 i_0_0_291 (.A1(poolingWindowX[16]), .A2(poolingWindowX[15]), .A3(
      poolingWindowX[14]), .A4(poolingWindowX[13]), .ZN(n_0_0_149));
   NOR4_X1 i_0_0_292 (.A1(poolingWindowX[12]), .A2(poolingWindowX[11]), .A3(
      poolingWindowX[10]), .A4(poolingWindowX[9]), .ZN(n_0_0_150));
   NAND2_X1 i_0_0_293 (.A1(n_0_0_153), .A2(n_0_0_152), .ZN(n_0_0_151));
   NOR4_X1 i_0_0_294 (.A1(poolingWindowX[24]), .A2(poolingWindowX[21]), .A3(
      poolingWindowX[19]), .A4(poolingWindowX[18]), .ZN(n_0_0_152));
   NOR2_X1 i_0_0_295 (.A1(poolingWindowX[27]), .A2(poolingWindowX[26]), .ZN(
      n_0_0_153));
   NAND3_X1 i_0_0_296 (.A1(n_0_0_157), .A2(n_0_0_156), .A3(n_0_0_155), .ZN(
      n_0_0_154));
   NOR4_X1 i_0_0_297 (.A1(poolingWindowX[23]), .A2(poolingWindowX[22]), .A3(
      poolingWindowX[20]), .A4(poolingWindowX[17]), .ZN(n_0_0_155));
   NOR2_X1 i_0_0_298 (.A1(poolingWindowX[28]), .A2(poolingWindowX[25]), .ZN(
      n_0_0_156));
   NOR2_X1 i_0_0_299 (.A1(poolingWindowX[30]), .A2(poolingWindowX[29]), .ZN(
      n_0_0_157));
   OAI21_X1 i_0_0_300 (.A(n_0_0_213), .B1(n_0_0_159), .B2(poolingWindowX[4]), 
      .ZN(n_0_0_158));
   AOI221_X1 i_0_0_301 (.A(n_0_0_160), .B1(n_0_0_161), .B2(n_0_0_214), .C1(
      n_0_0_228), .C2(n_0_0_162), .ZN(n_0_0_159));
   NOR3_X1 i_0_0_302 (.A1(n_0_0_30), .A2(poolingWindowX[2]), .A3(
      poolingWindowX[3]), .ZN(n_0_0_160));
   NAND2_X1 i_0_0_303 (.A1(poolingWindowX[2]), .A2(poolingWindowX[1]), .ZN(
      n_0_0_161));
   OAI21_X1 i_0_0_304 (.A(poolingWindowX[3]), .B1(poolingWindowX[2]), .B2(
      poolingWindowX[1]), .ZN(n_0_0_162));
   INV_X1 i_0_0_305 (.A(n_0_0_164), .ZN(n_0_0_163));
   NAND2_X1 i_0_0_306 (.A1(n_0_0_225), .A2(n_0_0_165), .ZN(n_0_0_164));
   NAND4_X1 i_0_0_307 (.A1(n_0_0_178), .A2(n_0_0_171), .A3(n_0_0_170), .A4(
      n_0_0_166), .ZN(n_0_0_165));
   NOR2_X1 i_0_0_308 (.A1(n_0_0_174), .A2(n_0_0_167), .ZN(n_0_0_166));
   NAND4_X1 i_0_0_309 (.A1(n_0_0_173), .A2(n_0_0_172), .A3(n_0_0_169), .A4(
      n_0_0_168), .ZN(n_0_0_167));
   NOR4_X1 i_0_0_310 (.A1(poolingWindowY[24]), .A2(poolingWindowY[21]), .A3(
      poolingWindowY[19]), .A4(poolingWindowY[18]), .ZN(n_0_0_168));
   NOR2_X1 i_0_0_311 (.A1(poolingWindowY[27]), .A2(poolingWindowY[26]), .ZN(
      n_0_0_169));
   NOR4_X1 i_0_0_312 (.A1(poolingWindowY[23]), .A2(poolingWindowY[22]), .A3(
      poolingWindowY[20]), .A4(poolingWindowY[17]), .ZN(n_0_0_170));
   NOR4_X1 i_0_0_313 (.A1(poolingWindowY[30]), .A2(poolingWindowY[29]), .A3(
      poolingWindowY[28]), .A4(poolingWindowY[25]), .ZN(n_0_0_171));
   NOR4_X1 i_0_0_314 (.A1(poolingWindowY[16]), .A2(poolingWindowY[15]), .A3(
      poolingWindowY[14]), .A4(poolingWindowY[13]), .ZN(n_0_0_172));
   NOR4_X1 i_0_0_315 (.A1(poolingWindowY[12]), .A2(poolingWindowY[11]), .A3(
      poolingWindowY[10]), .A4(poolingWindowY[9]), .ZN(n_0_0_173));
   NAND3_X1 i_0_0_316 (.A1(n_0_0_177), .A2(n_0_0_176), .A3(n_0_0_175), .ZN(
      n_0_0_174));
   NOR2_X1 i_0_0_317 (.A1(poolingWindowY[8]), .A2(poolingWindowY[5]), .ZN(
      n_0_0_175));
   NOR2_X1 i_0_0_318 (.A1(poolingWindowY[7]), .A2(poolingWindowY[6]), .ZN(
      n_0_0_176));
   NAND2_X1 i_0_0_319 (.A1(layerCounter[2]), .A2(n_0_0_28), .ZN(n_0_0_177));
   OAI21_X1 i_0_0_320 (.A(n_0_0_213), .B1(n_0_0_179), .B2(poolingWindowY[4]), 
      .ZN(n_0_0_178));
   AOI221_X1 i_0_0_321 (.A(n_0_0_180), .B1(n_0_0_181), .B2(n_0_0_214), .C1(
      n_0_0_228), .C2(n_0_0_182), .ZN(n_0_0_179));
   NOR3_X1 i_0_0_322 (.A1(n_0_0_30), .A2(poolingWindowY[2]), .A3(
      poolingWindowY[3]), .ZN(n_0_0_180));
   NAND2_X1 i_0_0_323 (.A1(poolingWindowY[2]), .A2(poolingWindowY[1]), .ZN(
      n_0_0_181));
   OAI21_X1 i_0_0_324 (.A(poolingWindowY[3]), .B1(poolingWindowY[2]), .B2(
      poolingWindowY[1]), .ZN(n_0_0_182));
   AOI21_X1 i_0_0_325 (.A(n_0_0_185), .B1(n_0_0_1), .B2(n_0_0_229), .ZN(
      n_0_0_183));
   OAI21_X1 i_0_0_326 (.A(n_0_0_221), .B1(n_0_0_185), .B2(n_0_0_184), .ZN(
      n_0_181));
   NAND2_X1 i_0_0_327 (.A1(n_0_0_229), .A2(n_0_0_1), .ZN(n_0_0_184));
   NAND2_X1 i_0_0_328 (.A1(n_0_0_222), .A2(start), .ZN(n_0_0_185));
   INV_X1 i_0_0_329 (.A(n_0_0_186), .ZN(n_0_143));
   NAND2_X1 i_0_0_330 (.A1(poolingReset), .A2(readAdress[0]), .ZN(n_0_0_186));
   INV_X1 i_0_0_331 (.A(n_0_0_187), .ZN(n_0_144));
   AOI21_X1 i_0_0_332 (.A(n_0_0_188), .B1(readAdress[1]), .B2(poolingReset), 
      .ZN(n_0_0_187));
   AOI21_X1 i_0_0_333 (.A(poolingReset), .B1(n_0_0_214), .B2(layerCounter[1]), 
      .ZN(n_0_0_188));
   NAND2_X1 i_0_0_334 (.A1(n_0_0_189), .A2(n_0_0_190), .ZN(n_0_145));
   AOI21_X1 i_0_0_335 (.A(n_0_0_191), .B1(readAdress[2]), .B2(poolingReset), 
      .ZN(n_0_0_189));
   NAND2_X1 i_0_0_336 (.A1(layerCounter[1]), .A2(n_0_0_200), .ZN(n_0_0_190));
   NOR3_X1 i_0_0_337 (.A1(n_0_0_196), .A2(poolingReset), .A3(layerCounter[2]), 
      .ZN(n_0_0_191));
   INV_X1 i_0_0_338 (.A(n_0_0_192), .ZN(n_0_162));
   AOI21_X1 i_0_0_339 (.A(n_0_0_199), .B1(readAdress[3]), .B2(poolingReset), 
      .ZN(n_0_0_192));
   NAND2_X1 i_0_0_340 (.A1(n_0_0_195), .A2(n_0_0_193), .ZN(n_0_163));
   NAND2_X1 i_0_0_341 (.A1(poolingReset), .A2(readAdress[4]), .ZN(n_0_0_193));
   NAND2_X1 i_0_0_342 (.A1(n_0_0_195), .A2(n_0_0_194), .ZN(n_0_164));
   NAND2_X1 i_0_0_343 (.A1(poolingReset), .A2(readAdress[5]), .ZN(n_0_0_194));
   NAND2_X1 i_0_0_344 (.A1(n_0_0_199), .A2(n_0_0_27), .ZN(n_0_0_195));
   NAND3_X1 i_0_0_345 (.A1(n_0_0_227), .A2(layerCounter[0]), .A3(layerCounter[2]), 
      .ZN(n_0_0_27));
   NAND2_X1 i_0_0_346 (.A1(n_0_0_227), .A2(layerCounter[0]), .ZN(n_0_0_196));
   OAI21_X1 i_0_0_347 (.A(n_0_0_197), .B1(n_0_0_31), .B2(poolingReset), .ZN(
      n_0_165));
   NAND2_X1 i_0_0_348 (.A1(poolingReset), .A2(readAdress[6]), .ZN(n_0_0_197));
   OAI21_X1 i_0_0_349 (.A(n_0_0_198), .B1(n_0_0_31), .B2(poolingReset), .ZN(
      n_0_166));
   NAND2_X1 i_0_0_350 (.A1(poolingReset), .A2(readAdress[7]), .ZN(n_0_0_198));
   MUX2_X1 i_0_0_351 (.A(n_0_0_36), .B(readAdress[8]), .S(poolingReset), 
      .Z(n_0_167));
   NOR2_X1 i_0_0_352 (.A1(n_0_0_202), .A2(n_0_0_201), .ZN(n_0_168));
   NOR2_X1 i_0_0_353 (.A1(poolingReset), .A2(n_0_178), .ZN(n_0_0_199));
   NOR2_X1 i_0_0_354 (.A1(n_0_0_228), .A2(poolingReset), .ZN(n_0_0_200));
   NOR3_X1 i_0_0_355 (.A1(n_0_0_213), .A2(n_0_0_0), .A3(poolingReset), .ZN(
      n_0_0_201));
   AOI21_X1 i_0_0_356 (.A(n_0_0_204), .B1(readAdress[9]), .B2(poolingReset), 
      .ZN(n_0_0_202));
   INV_X1 i_0_0_357 (.A(n_0_0_203), .ZN(n_0_169));
   AOI21_X1 i_0_0_358 (.A(n_0_0_204), .B1(readAdress[10]), .B2(poolingReset), 
      .ZN(n_0_0_203));
   NOR2_X1 i_0_0_359 (.A1(poolingReset), .A2(n_0_0_25), .ZN(n_0_0_204));
   AND2_X1 i_0_0_360 (.A1(n_0_0_213), .A2(n_0_0_0), .ZN(n_0_0_25));
   MUX2_X1 i_0_0_361 (.A(n_0_0_37), .B(readAdress[11]), .S(poolingReset), 
      .Z(n_0_170));
   MUX2_X1 i_0_0_362 (.A(n_0_0_38), .B(readAdress[12]), .S(poolingReset), 
      .Z(n_0_171));
   MUX2_X1 i_0_0_363 (.A(n_0_0_39), .B(readAdress[13]), .S(poolingReset), 
      .Z(n_0_172));
   INV_X1 i_0_0_364 (.A(n_0_0_205), .ZN(n_0_173));
   AOI21_X1 i_0_0_365 (.A(n_0_0_207), .B1(readAdress[14]), .B2(poolingReset), 
      .ZN(n_0_0_205));
   INV_X1 i_0_0_366 (.A(n_0_0_206), .ZN(n_0_174));
   AOI21_X1 i_0_0_367 (.A(n_0_0_207), .B1(readAdress[15]), .B2(poolingReset), 
      .ZN(n_0_0_206));
   NOR2_X1 i_0_0_368 (.A1(poolingReset), .A2(n_0_0_208), .ZN(n_0_0_207));
   XOR2_X1 i_0_0_369 (.A(n_0_0_4), .B(n_0_0_209), .Z(n_0_0_208));
   NAND2_X1 i_0_0_370 (.A1(n_0_0_30), .A2(n_0_0_26), .ZN(n_0_0_209));
   NAND2_X1 i_0_0_371 (.A1(n_0_0_28), .A2(n_0_0_228), .ZN(n_0_0_26));
   NOR2_X1 i_0_0_372 (.A1(n_0_0_28), .A2(n_0_0_228), .ZN(n_0_175));
   NOR2_X1 i_0_0_373 (.A1(n_0_0_227), .A2(n_0_0_226), .ZN(n_0_0_28));
   NAND2_X1 i_0_0_374 (.A1(n_0_0_29), .A2(n_0_0_210), .ZN(n_0_176));
   NAND2_X1 i_0_0_375 (.A1(layerCounter[1]), .A2(n_0_0_214), .ZN(n_0_0_210));
   NAND2_X1 i_0_0_376 (.A1(n_0_0_228), .A2(layerCounter[1]), .ZN(n_0_0_211));
   NAND2_X1 i_0_0_377 (.A1(n_0_0_226), .A2(layerCounter[1]), .ZN(n_0_0_212));
   NAND2_X1 i_0_0_378 (.A1(layerCounter[2]), .A2(n_0_0_31), .ZN(n_0_0_29));
   NOR2_X1 i_0_0_379 (.A1(layerCounter[2]), .A2(n_0_0_31), .ZN(n_0_177));
   INV_X1 i_0_0_380 (.A(n_0_0_213), .ZN(n_0_178));
   NAND2_X1 i_0_0_381 (.A1(n_0_0_31), .A2(n_0_0_228), .ZN(n_0_0_213));
   NOR2_X1 i_0_0_382 (.A1(layerCounter[2]), .A2(layerCounter[0]), .ZN(n_0_0_214));
   INV_X1 i_0_0_383 (.A(n_0_0_31), .ZN(n_0_0_30));
   NOR2_X1 i_0_0_384 (.A1(layerCounter[1]), .A2(layerCounter[0]), .ZN(n_0_0_31));
   INV_X1 i_0_0_385 (.A(n_0_0_43), .ZN(n_0_0_215));
   INV_X1 i_0_0_386 (.A(n_0_0_42), .ZN(n_0_0_216));
   INV_X1 i_0_0_387 (.A(writeAdress[1]), .ZN(n_0_0_217));
   INV_X1 i_0_0_388 (.A(writeAdress[3]), .ZN(n_0_0_218));
   INV_X1 i_0_0_389 (.A(writeAdress[4]), .ZN(n_0_0_219));
   INV_X1 i_0_0_390 (.A(writeAdress[5]), .ZN(n_0_0_220));
   INV_X1 i_0_0_391 (.A(reset), .ZN(n_0_0_221));
   INV_X1 i_0_0_392 (.A(DMA_start), .ZN(n_0_0_222));
   INV_X1 i_0_0_393 (.A(poolingState[0]), .ZN(n_0_0_223));
   INV_X1 i_0_0_394 (.A(poolingCounter[0]), .ZN(n_0_0_224));
   INV_X1 i_0_0_395 (.A(poolingWindowY[31]), .ZN(n_0_0_225));
   INV_X1 i_0_0_396 (.A(layerCounter[0]), .ZN(n_0_0_226));
   INV_X1 i_0_0_397 (.A(layerCounter[1]), .ZN(n_0_0_227));
   INV_X1 i_0_0_398 (.A(layerCounter[2]), .ZN(n_0_0_228));
   INV_X1 i_0_0_399 (.A(layerCounter[31]), .ZN(n_0_0_229));
   NOR2_X1 i_0_0_400 (.A1(n_0_0_186), .A2(poolingState[0]), .ZN(n_0_201));
   CLKGATETST_X1 clk_gate_DMA_offset_reg (.CK(clk), .E(n_0_139), .SE(1'b0), 
      .GCK(n_0_179));
   MUX2_X1 finishCNN_reg_enable_mux_0 (.A(finish), .B(n_0_36), .S(n_0_181), 
      .Z(n_0_182));
   MUX2_X1 DMA_start_reg_enable_mux_0 (.A(DMA_start), .B(n_0_37), .S(n_0_180), 
      .Z(n_0_199));
   MUX2_X1 \poolingState_reg[0]_enable_mux_0  (.A(poolingState[0]), .B(n_0_38), 
      .S(n_0_142), .Z(n_0_200));
   MUX2_X1 poolingReset_reg_enable_mux_0 (.A(poolingReset), .B(n_0_140), 
      .S(n_0_141), .Z(n_0_217));
endmodule
