
// 	Wed May  5 21:37:16 2021
//	vlsi
//	localhost.localdomain

module Booth_Multiplier (multiplicand, multiplier, product);

output [15:0] product;
input [7:0] multiplicand;
input [7:0] multiplier;
wire n_0_0_77;
wire n_0_0_2;
wire n_0_0_78;
wire n_0_0_3;
wire n_0_0_79;
wire n_0_0_4;
wire n_0_0_80;
wire n_0_0_5;
wire n_0_0_81;
wire n_0_0_6;
wire n_0_0_82;
wire n_0_0_0;
wire n_0_0_83;
wire n_0_0_1;
wire n_0_0_84;
wire n_0_0_7;
wire n_0_0_85;
wire n_0_0_8;
wire n_0_0_86;
wire n_0_0_9;
wire n_0_0_87;
wire n_0_0_10;
wire n_0_0_88;
wire n_0_0_11;
wire n_0_0_89;
wire n_0_0_12;
wire n_0_0_90;
wire n_0_0_13;
wire n_0_0_91;
wire n_0_0_14;
wire n_0_0_92;
wire n_0_0_15;
wire n_0_0_93;
wire n_0_0_16;
wire n_0_0_94;
wire n_0_0_17;
wire n_0_0_95;
wire n_0_0_18;
wire n_0_0_96;
wire n_0_0_19;
wire n_0_0_97;
wire n_0_0_20;
wire n_0_0_98;
wire n_0_0_21;
wire n_0_0_99;
wire n_0_0_22;
wire n_0_0_100;
wire n_0_0_23;
wire n_0_0_101;
wire n_0_0_24;
wire n_0_0_102;
wire n_0_0_25;
wire n_0_0_103;
wire n_0_0_26;
wire n_0_0_104;
wire n_0_0_27;
wire n_0_0_105;
wire n_0_0_28;
wire n_0_0_106;
wire n_0_0_29;
wire n_0_0_107;
wire n_0_0_30;
wire n_0_0_108;
wire n_0_0_31;
wire n_0_0_109;
wire n_0_0_32;
wire n_0_0_110;
wire n_0_0_33;
wire n_0_0_111;
wire n_0_0_34;
wire n_0_0_112;
wire n_0_0_35;
wire n_0_0_113;
wire n_0_0_36;
wire n_0_0_114;
wire n_0_0_37;
wire n_0_0_115;
wire n_0_0_38;
wire n_0_0_116;
wire n_0_0_39;
wire n_0_0_117;
wire n_0_0_40;
wire n_0_0_118;
wire n_0_0_41;
wire n_0_0_119;
wire n_0_0_42;
wire n_0_0_120;
wire n_0_0_43;
wire n_0_0_121;
wire n_0_0_44;
wire n_0_0_122;
wire n_0_0_45;
wire n_0_0_123;
wire n_0_0_46;
wire n_0_0_124;
wire n_0_0_47;
wire n_0_0_125;
wire n_0_0_48;
wire n_0_0_126;
wire n_0_0_49;
wire n_0_0_127;
wire n_0_0_50;
wire n_0_0_128;
wire n_0_0_51;
wire n_0_0_129;
wire n_0_0_52;
wire n_0_0_130;
wire n_0_0_53;
wire n_0_0_131;
wire n_0_0_54;
wire n_0_0_132;
wire n_0_0_55;
wire n_0_0_133;
wire n_0_0_56;
wire n_0_0_134;
wire n_0_0_57;
wire n_0_0_135;
wire n_0_0_58;
wire n_0_0_136;
wire n_0_0_59;
wire n_0_0_137;
wire n_0_0_60;
wire n_0_0_138;
wire n_0_0_61;
wire n_0_0_139;
wire n_0_0_62;
wire n_0_0_140;
wire n_0_0_63;
wire n_0_0_141;
wire n_0_0_64;
wire n_0_0_142;
wire n_0_0_65;
wire n_0_0_143;
wire n_0_0_66;
wire n_0_0_144;
wire n_0_0_67;
wire n_0_0_145;
wire n_0_0_68;
wire n_0_0_146;
wire n_0_0_69;
wire n_0_0_147;
wire n_0_0_70;
wire n_0_0_148;
wire n_0_0_71;
wire n_0_0_149;
wire n_0_0_72;
wire n_0_0_150;
wire n_0_0_73;
wire n_0_0_151;
wire n_0_0_74;
wire n_0_0_152;
wire n_0_0_75;
wire n_0_0_153;
wire n_0_0_76;
wire n_0_0_154;
wire n_0_0_155;
wire n_0_0_156;
wire n_0_0_157;
wire n_0_0_158;
wire n_0_0_159;
wire n_0_0_160;
wire n_0_0_161;
wire n_0_0_162;
wire n_0_0_163;
wire n_0_0_164;
wire n_0_0_165;
wire n_0_0_166;
wire n_0_0_167;
wire n_0_0_168;
wire n_0_0_169;
wire n_0_0_170;
wire n_0_0_171;
wire n_0_0_172;
wire n_0_0_173;
wire n_0_0_174;
wire n_0_0_175;
wire n_0_0_176;
wire n_0_0_177;
wire n_0_0_178;
wire n_0_0_179;
wire n_0_0_180;
wire n_0_0_181;
wire n_0_0_182;
wire n_0_0_183;
wire n_0_0_184;
wire n_0_0_185;
wire n_0_0_186;
wire n_0_0_187;
wire n_0_0_188;
wire n_0_0_189;
wire n_0_0_190;
wire n_0_0_191;
wire n_0_0_192;
wire n_0_0_193;
wire n_0_0_194;
wire n_0_0_195;
wire n_0_0_196;
wire n_0_0_197;
wire n_0_0_198;
wire n_0_0_199;
wire n_0_0_200;
wire n_0_0_201;
wire n_0_0_202;
wire n_0_0_203;
wire n_0_0_204;
wire n_0_0_205;
wire n_0_0_206;
wire n_0_0_207;
wire n_0_0_208;
wire n_0_0_209;
wire n_0_0_210;
wire n_0_0_211;
wire n_0_0_212;
wire n_0_0_213;
wire n_0_0_214;
wire n_0_0_215;
wire n_0_0_216;
wire n_0_0_217;
wire n_0_0_218;
wire n_0_0_219;
wire n_0_0_220;
wire n_0_0_221;
wire n_0_0_222;
wire n_0_0_223;
wire n_0_0_224;
wire n_0_0_225;
wire n_0_0_226;
wire n_0_0_227;
wire n_0_0_228;
wire n_0_0_229;
wire n_0_0_230;
wire n_0_0_231;
wire n_0_0_232;
wire n_0_0_233;
wire n_0_0_234;
wire n_0_0_235;
wire n_0_0_236;
wire n_0_0_237;
wire n_0_0_238;
wire n_0_0_239;
wire n_0_0_240;
wire n_0_0_241;
wire n_0_0_242;
wire n_0_0_243;
wire n_0_0_244;
wire n_0_0_245;
wire n_0_0_246;
wire n_0_0_247;
wire n_0_0_248;
wire n_0_0_249;
wire n_0_0_250;
wire n_0_0_251;
wire n_0_0_252;
wire n_0_0_253;
wire n_0_0_254;
wire n_0_0_255;
wire n_0_0_256;
wire n_0_0_257;
wire n_0_0_258;
wire n_0_0_259;
wire n_0_0_260;
wire n_0_0_261;
wire n_0_0_262;
wire n_0_0_263;
wire n_0_0_264;
wire n_0_0_265;
wire n_0_0_266;
wire n_0_0_267;
wire n_0_0_268;
wire n_0_0_269;
wire n_0_0_270;
wire n_0_0_271;
wire n_0_0_272;
wire n_0_0_273;
wire n_0_0_274;
wire n_0_0_275;
wire n_0_0_276;
wire n_0_0_277;
wire n_0_0_278;
wire n_0_0_279;
wire n_0_0_280;
wire n_0_0_281;
wire n_0_0_282;
wire n_0_0_283;
wire n_0_0_284;
wire n_0_0_285;
wire n_0_0_286;
wire n_0_0_287;
wire n_0_0_288;
wire n_0_0_289;
wire n_0_0_290;
wire n_0_0_291;
wire n_0_0_292;
wire n_0_0_293;
wire n_0_0_294;
wire n_0_0_295;
wire n_0_0_296;
wire n_0_0_297;
wire n_0_0_298;
wire n_0_0_299;
wire n_0_0_300;
wire n_0_0_301;
wire n_0_0_302;
wire n_0_0_303;
wire n_0_0_304;
wire n_0_0_305;
wire n_0_0_306;
wire n_0_0_307;
wire n_0_0_308;
wire n_0_0_309;
wire n_0_0_310;
wire n_0_0_311;
wire n_0_0_312;
wire n_0_0_313;
wire n_0_0_314;
wire n_0_0_315;
wire n_0_0_316;
wire n_0_0_317;
wire n_0_0_318;
wire n_0_0_319;
wire n_0_0_320;
wire n_0_0_321;
wire n_0_0_322;
wire n_0_0_323;
wire n_0_0_324;
wire n_0_0_325;
wire n_0_0_326;
wire n_0_0_327;
wire n_0_0_328;
wire n_0_0_329;
wire n_0_0_330;
wire n_0_0_331;
wire n_0_0_332;
wire n_0_0_333;
wire n_0_0_334;
wire n_0_0_335;
wire n_0_0_336;
wire n_0_0_337;
wire n_0_0_338;
wire n_0_0_339;
wire n_0_0_340;
wire n_0_0_341;
wire n_0_0_342;
wire n_0_0_343;
wire n_0_0_344;
wire n_0_0_345;
wire n_0_0_346;
wire n_0_0_347;
wire n_0_0_348;
wire n_0_0_349;
wire n_0_0_350;
wire n_0_0_351;
wire n_0_0_352;
wire n_0_0_353;
wire n_0_0_354;
wire n_0_0_355;
wire n_0_0_356;
wire n_0_0_357;
wire n_0_0_358;
wire n_0_0_359;
wire n_0_0_360;
wire n_0_0_361;
wire n_0_0_362;
wire n_0_0_363;
wire n_0_0_364;
wire n_0_0_365;
wire n_0_0_366;
wire n_0_0_367;
wire n_0_0_368;
wire n_0_0_369;
wire n_0_0_370;
wire n_0_0_371;
wire n_0_0_372;
wire n_0_0_373;
wire n_0_0_374;
wire n_0_0_375;
wire n_0_0_376;
wire n_0_0_377;
wire n_0_0_378;
wire n_0_0_379;
wire n_0_0_380;
wire n_0_0_381;
wire n_0_0_382;
wire n_0_0_383;
wire n_0_0_384;
wire n_0_0_385;
wire n_0_0_386;
wire n_0_0_387;
wire n_0_0_388;
wire n_0_0_389;
wire n_0_0_390;
wire n_0_0_391;
wire n_0_0_392;
wire n_0_0_393;
wire n_0_0_394;
wire spc__n1;
wire spc__n2;
wire spc__n3;
wire spc__n4;
wire spc__n5;
wire spc__n6;
wire spc__n7;
wire spc__n8;
wire spc__n9;
wire spt__n28;
wire spt__n31;
wire spt__n36;
wire spt__n41;
wire spw__n66;
wire spw__n69;
wire spw__n105;
wire spw__n162;
wire spw__n163;
wire spw__n164;
wire spw__n165;
wire spw__n166;
wire spw__n572;
wire spw__n573;
wire spw__n574;
wire spw__n575;
wire spw__n576;
wire spw__n577;
wire spw__n578;
wire spw__n579;
wire spw__n580;
wire spw__n581;
wire spw__n582;
wire spw__n583;
wire spw__n584;
wire spw__n662;
wire spw__n682;
wire spw__n683;
wire spw__n684;
wire spw__n685;
wire spw__n686;
wire spw__n687;
wire spw__n688;
wire spw__n689;
wire spw__n690;
wire spw__n691;
wire spw__n692;

// WARNING . Detected multiport output net(s). Introducing ASSIGN statements.
// This may cause simulation/synthesis mismatches . 
assign product[15] = product[14];

INV_X1 i_0_0_332 (.ZN (n_0_0_394), .A (multiplicand[6]));
INV_X1 i_0_0_331 (.ZN (n_0_0_393), .A (multiplier[6]));
INV_X1 i_0_0_330 (.ZN (n_0_0_392), .A (multiplier[5]));
INV_X1 i_0_0_329 (.ZN (n_0_0_391), .A (multiplier[4]));
INV_X1 i_0_0_328 (.ZN (n_0_0_390), .A (multiplier[3]));
INV_X1 i_0_0_327 (.ZN (n_0_0_389), .A (multiplier[2]));
INV_X1 i_0_0_326 (.ZN (n_0_0_388), .A (multiplier[1]));
INV_X1 i_0_0_325 (.ZN (n_0_0_387), .A (n_0_0_6));
INV_X1 i_0_0_324 (.ZN (n_0_0_386), .A (n_0_0_9));
INV_X1 i_0_0_323 (.ZN (n_0_0_385), .A (n_0_0_14));
INV_X1 i_0_0_322 (.ZN (n_0_0_384), .A (n_0_0_24));
INV_X1 i_0_0_321 (.ZN (n_0_0_383), .A (n_0_0_34));
INV_X1 i_0_0_320 (.ZN (n_0_0_382), .A (n_0_0_44));
INV_X1 i_0_0_319 (.ZN (n_0_0_381), .A (n_0_0_49));
INV_X1 i_0_0_318 (.ZN (n_0_0_380), .A (n_0_0_54));
INV_X1 i_0_0_317 (.ZN (n_0_0_379), .A (n_0_0_64));
INV_X1 i_0_0_316 (.ZN (n_0_0_378), .A (n_0_0_69));
NOR2_X4 i_0_0_315 (.ZN (n_0_0_377), .A1 (multiplicand[1]), .A2 (multiplicand[0]));
INV_X2 i_0_0_314 (.ZN (n_0_0_376), .A (n_0_0_377));
NOR2_X4 i_0_0_313 (.ZN (n_0_0_375), .A1 (multiplicand[2]), .A2 (n_0_0_376));
INV_X1 i_0_0_312 (.ZN (n_0_0_374), .A (n_0_0_375));
NOR2_X2 i_0_0_311 (.ZN (n_0_0_373), .A1 (multiplicand[3]), .A2 (n_0_0_374));
INV_X1 i_0_0_310 (.ZN (n_0_0_372), .A (n_0_0_373));
NOR2_X1 i_0_0_309 (.ZN (n_0_0_371), .A1 (multiplicand[4]), .A2 (n_0_0_372));
INV_X1 i_0_0_308 (.ZN (n_0_0_370), .A (n_0_0_371));
NOR2_X1 i_0_0_307 (.ZN (n_0_0_369), .A1 (multiplicand[5]), .A2 (n_0_0_370));
OAI21_X1 i_0_0_306 (.ZN (n_0_0_368), .A (multiplicand[6]), .B1 (multiplicand[5]), .B2 (n_0_0_370));
NAND2_X1 i_0_0_305 (.ZN (n_0_0_367), .A1 (n_0_0_394), .A2 (n_0_0_369));
NAND2_X4 i_0_0_304 (.ZN (n_0_0_366), .A1 (n_0_0_368), .A2 (n_0_0_367));
INV_X4 i_0_0_303 (.ZN (n_0_0_365), .A (n_0_0_366));
XNOR2_X1 i_0_0_302 (.ZN (n_0_0_364), .A (multiplicand[7]), .B (n_0_0_368));
INV_X1 i_0_0_301 (.ZN (n_0_0_363), .A (n_0_0_364));
NAND2_X1 i_0_0_300 (.ZN (n_0_0_362), .A1 (multiplier[5]), .A2 (n_0_0_391));
INV_X1 i_0_0_299 (.ZN (n_0_0_361), .A (n_0_0_362));
NAND2_X1 i_0_0_298 (.ZN (n_0_0_360), .A1 (multiplier[4]), .A2 (n_0_0_390));
INV_X1 i_0_0_297 (.ZN (n_0_0_359), .A (n_0_0_360));
NAND2_X1 i_0_0_296 (.ZN (n_0_0_358), .A1 (multiplier[3]), .A2 (n_0_0_389));
INV_X1 i_0_0_295 (.ZN (n_0_0_357), .A (n_0_0_358));
OAI21_X1 i_0_0_294 (.ZN (n_0_0_356), .A (multiplier[0]), .B1 (multiplicand[7]), .B2 (n_0_0_367));
AOI21_X1 i_0_0_293 (.ZN (n_0_0_355), .A (n_0_0_356), .B1 (multiplicand[7]), .B2 (n_0_0_367));
INV_X1 i_0_0_292 (.ZN (n_0_0_354), .A (n_0_0_355));
NAND2_X1 i_0_0_291 (.ZN (n_0_0_353), .A1 (multiplicand[6]), .A2 (n_0_0_354));
NAND2_X1 i_0_0_290 (.ZN (n_0_0_352), .A1 (n_0_0_394), .A2 (n_0_0_355));
OAI22_X1 i_0_0_289 (.ZN (n_0_0_351), .A1 (n_0_0_386), .A2 (n_0_0_353), .B1 (n_0_0_9), .B2 (n_0_0_352));
AND2_X1 i_0_0_288 (.ZN (n_0_0_350), .A1 (n_0_0_388), .A2 (multiplier[0]));
XOR2_X1 i_0_0_287 (.Z (n_0_0_349), .A (multiplicand[7]), .B (n_0_0_351));
NOR2_X1 i_0_0_286 (.ZN (n_0_0_348), .A1 (n_0_0_388), .A2 (n_0_0_354));
AOI21_X1 i_0_0_285 (.ZN (n_0_0_347), .A (n_0_0_355), .B1 (n_0_0_387), .B2 (n_0_0_365));
AOI21_X1 i_0_0_284 (.ZN (n_0_0_346), .A (n_0_0_347), .B1 (n_0_0_6), .B2 (n_0_0_366));
NOR2_X1 i_0_0_283 (.ZN (n_0_0_345), .A1 (n_0_0_388), .A2 (multiplier[0]));
XNOR2_X1 i_0_0_282 (.ZN (n_0_0_344), .A (n_0_0_363), .B (n_0_0_346));
AOI221_X1 i_0_0_281 (.ZN (n_0_0_343), .A (n_0_0_348), .B1 (n_0_0_345), .B2 (n_0_0_344)
    , .C1 (n_0_0_350), .C2 (n_0_0_349));
INV_X1 i_0_0_280 (.ZN (n_0_0_342), .A (n_0_0_343));
NOR2_X1 i_0_0_279 (.ZN (n_0_0_341), .A1 (multiplicand[6]), .A2 (n_0_0_19));
AND2_X2 i_0_0_278 (.ZN (n_0_0_340), .A1 (multiplicand[6]), .A2 (n_0_0_19));
OAI22_X1 i_0_0_277 (.ZN (n_0_0_339), .A1 (n_0_0_343), .A2 (n_0_0_341), .B1 (n_0_0_342), .B2 (n_0_0_340));
NAND2_X1 i_0_0_276 (.ZN (n_0_0_338), .A1 (n_0_0_389), .A2 (multiplier[1]));
INV_X1 i_0_0_275 (.ZN (n_0_0_337), .A (n_0_0_338));
XNOR2_X1 i_0_0_274 (.ZN (n_0_0_336), .A (multiplicand[7]), .B (n_0_0_339));
NAND2_X1 i_0_0_273 (.ZN (n_0_0_335), .A1 (multiplier[2]), .A2 (n_0_0_388));
INV_X1 i_0_0_272 (.ZN (n_0_0_334), .A (n_0_0_335));
NAND2_X1 i_0_0_271 (.ZN (n_0_0_333), .A1 (n_0_0_338), .A2 (n_0_0_335));
AOI21_X1 i_0_0_270 (.ZN (n_0_0_332), .A (n_0_0_342), .B1 (n_0_0_385), .B2 (n_0_0_365));
AOI21_X1 i_0_0_269 (.ZN (n_0_0_331), .A (n_0_0_332), .B1 (n_0_0_14), .B2 (n_0_0_366));
XOR2_X1 i_0_0_268 (.Z (n_0_0_330), .A (n_0_0_364), .B (n_0_0_331));
AOI22_X1 i_0_0_267 (.ZN (n_0_0_329), .A1 (n_0_0_337), .A2 (n_0_0_336), .B1 (n_0_0_334), .B2 (n_0_0_330));
OAI21_X1 i_0_0_266 (.ZN (n_0_0_328), .A (n_0_0_329), .B1 (n_0_0_343), .B2 (n_0_0_333));
INV_X1 i_0_0_265 (.ZN (n_0_0_327), .A (n_0_0_328));
AOI21_X1 i_0_0_264 (.ZN (n_0_0_326), .A (n_0_0_327), .B1 (n_0_0_24), .B2 (n_0_0_366));
AOI21_X1 i_0_0_263 (.ZN (n_0_0_325), .A (n_0_0_326), .B1 (n_0_0_384), .B2 (n_0_0_365));
XOR2_X1 i_0_0_262 (.Z (n_0_0_324), .A (n_0_0_363), .B (n_0_0_325));
NOR2_X1 i_0_0_261 (.ZN (n_0_0_323), .A1 (multiplicand[6]), .A2 (n_0_0_29));
AND2_X1 i_0_0_260 (.ZN (n_0_0_322), .A1 (multiplicand[6]), .A2 (n_0_0_29));
OAI22_X1 i_0_0_259 (.ZN (n_0_0_321), .A1 (n_0_0_327), .A2 (n_0_0_323), .B1 (n_0_0_328), .B2 (n_0_0_322));
NAND2_X1 i_0_0_258 (.ZN (n_0_0_320), .A1 (n_0_0_390), .A2 (multiplier[2]));
INV_X1 i_0_0_257 (.ZN (n_0_0_319), .A (n_0_0_320));
XNOR2_X1 i_0_0_256 (.ZN (n_0_0_318), .A (multiplicand[7]), .B (n_0_0_321));
NAND2_X1 i_0_0_255 (.ZN (n_0_0_317), .A1 (n_0_0_358), .A2 (n_0_0_320));
INV_X1 i_0_0_254 (.ZN (n_0_0_316), .A (n_0_0_317));
AOI222_X1 i_0_0_253 (.ZN (n_0_0_315), .A1 (n_0_0_319), .A2 (n_0_0_318), .B1 (n_0_0_328)
    , .B2 (n_0_0_316), .C1 (n_0_0_357), .C2 (n_0_0_324));
INV_X1 i_0_0_252 (.ZN (n_0_0_314), .A (n_0_0_315));
AOI21_X1 i_0_0_251 (.ZN (n_0_0_313), .A (n_0_0_315), .B1 (n_0_0_34), .B2 (n_0_0_366));
AOI21_X1 i_0_0_250 (.ZN (n_0_0_312), .A (n_0_0_313), .B1 (n_0_0_383), .B2 (n_0_0_365));
XOR2_X1 i_0_0_249 (.Z (n_0_0_311), .A (n_0_0_363), .B (n_0_0_312));
NAND2_X1 i_0_0_248 (.ZN (n_0_0_310), .A1 (n_0_0_391), .A2 (multiplier[3]));
INV_X1 i_0_0_247 (.ZN (n_0_0_309), .A (n_0_0_310));
NAND2_X1 i_0_0_246 (.ZN (n_0_0_308), .A1 (n_0_0_360), .A2 (n_0_0_310));
INV_X1 i_0_0_245 (.ZN (n_0_0_307), .A (n_0_0_308));
NOR2_X1 i_0_0_244 (.ZN (n_0_0_306), .A1 (multiplicand[6]), .A2 (n_0_0_39));
AND2_X2 i_0_0_243 (.ZN (n_0_0_305), .A1 (multiplicand[6]), .A2 (n_0_0_39));
OAI22_X1 i_0_0_242 (.ZN (n_0_0_304), .A1 (n_0_0_315), .A2 (n_0_0_306), .B1 (n_0_0_314), .B2 (n_0_0_305));
XNOR2_X1 i_0_0_241 (.ZN (n_0_0_303), .A (multiplicand[7]), .B (n_0_0_304));
AOI222_X1 i_0_0_240 (.ZN (n_0_0_302), .A1 (n_0_0_314), .A2 (n_0_0_307), .B1 (n_0_0_309)
    , .B2 (n_0_0_303), .C1 (n_0_0_359), .C2 (n_0_0_311));
INV_X1 i_0_0_239 (.ZN (n_0_0_301), .A (n_0_0_302));
AOI21_X1 i_0_0_238 (.ZN (n_0_0_300), .A (n_0_0_302), .B1 (n_0_0_44), .B2 (n_0_0_366));
AOI21_X1 i_0_0_237 (.ZN (n_0_0_299), .A (n_0_0_300), .B1 (n_0_0_382), .B2 (n_0_0_365));
XOR2_X1 i_0_0_236 (.Z (n_0_0_298), .A (n_0_0_363), .B (n_0_0_299));
OAI33_X1 i_0_0_235 (.ZN (n_0_0_297), .A1 (n_0_0_394), .A2 (n_0_0_381), .A3 (n_0_0_301)
    , .B1 (multiplicand[6]), .B2 (n_0_0_49), .B3 (n_0_0_302));
NAND2_X1 i_0_0_234 (.ZN (n_0_0_296), .A1 (n_0_0_392), .A2 (multiplier[4]));
INV_X1 i_0_0_233 (.ZN (n_0_0_295), .A (n_0_0_296));
XOR2_X1 i_0_0_232 (.Z (n_0_0_294), .A (multiplicand[7]), .B (n_0_0_297));
NAND2_X1 i_0_0_231 (.ZN (n_0_0_293), .A1 (n_0_0_362), .A2 (n_0_0_296));
INV_X1 i_0_0_230 (.ZN (n_0_0_292), .A (n_0_0_293));
AOI222_X1 i_0_0_229 (.ZN (n_0_0_291), .A1 (n_0_0_295), .A2 (n_0_0_294), .B1 (n_0_0_301)
    , .B2 (n_0_0_292), .C1 (n_0_0_361), .C2 (n_0_0_298));
INV_X1 i_0_0_228 (.ZN (n_0_0_290), .A (n_0_0_291));
AOI21_X1 i_0_0_227 (.ZN (n_0_0_289), .A (n_0_0_290), .B1 (n_0_0_380), .B2 (n_0_0_365));
AOI21_X1 i_0_0_226 (.ZN (n_0_0_288), .A (n_0_0_289), .B1 (n_0_0_54), .B2 (n_0_0_366));
NAND2_X1 i_0_0_225 (.ZN (n_0_0_287), .A1 (multiplier[6]), .A2 (n_0_0_392));
INV_X1 i_0_0_224 (.ZN (n_0_0_286), .A (n_0_0_287));
XOR2_X1 i_0_0_223 (.Z (n_0_0_285), .A (n_0_0_364), .B (n_0_0_288));
NOR2_X1 i_0_0_222 (.ZN (n_0_0_284), .A1 (multiplicand[6]), .A2 (n_0_0_59));
AND2_X1 i_0_0_221 (.ZN (n_0_0_283), .A1 (multiplicand[6]), .A2 (n_0_0_59));
OAI22_X1 i_0_0_220 (.ZN (n_0_0_282), .A1 (n_0_0_291), .A2 (n_0_0_284), .B1 (n_0_0_290), .B2 (n_0_0_283));
NAND2_X1 i_0_0_219 (.ZN (n_0_0_281), .A1 (n_0_0_393), .A2 (multiplier[5]));
INV_X1 i_0_0_218 (.ZN (n_0_0_280), .A (n_0_0_281));
XNOR2_X1 i_0_0_217 (.ZN (n_0_0_279), .A (multiplicand[7]), .B (n_0_0_282));
NAND2_X1 i_0_0_216 (.ZN (n_0_0_278), .A1 (n_0_0_287), .A2 (n_0_0_281));
INV_X1 i_0_0_215 (.ZN (n_0_0_277), .A (n_0_0_278));
AOI222_X1 i_0_0_214 (.ZN (n_0_0_276), .A1 (n_0_0_280), .A2 (n_0_0_279), .B1 (n_0_0_290)
    , .B2 (n_0_0_277), .C1 (n_0_0_286), .C2 (n_0_0_285));
INV_X1 i_0_0_213 (.ZN (n_0_0_275), .A (n_0_0_276));
OAI33_X1 i_0_0_212 (.ZN (n_0_0_274), .A1 (n_0_0_394), .A2 (n_0_0_378), .A3 (n_0_0_275)
    , .B1 (multiplicand[6]), .B2 (n_0_0_69), .B3 (n_0_0_276));
NOR2_X1 i_0_0_211 (.ZN (n_0_0_273), .A1 (multiplier[7]), .A2 (n_0_0_393));
INV_X1 i_0_0_210 (.ZN (n_0_0_272), .A (n_0_0_273));
XOR2_X1 i_0_0_209 (.Z (n_0_0_271), .A (multiplicand[7]), .B (n_0_0_274));
NAND2_X1 i_0_0_208 (.ZN (n_0_0_270), .A1 (multiplier[7]), .A2 (n_0_0_393));
INV_X1 i_0_0_207 (.ZN (n_0_0_269), .A (n_0_0_270));
NAND2_X1 i_0_0_206 (.ZN (n_0_0_268), .A1 (n_0_0_272), .A2 (n_0_0_270));
INV_X1 i_0_0_205 (.ZN (n_0_0_267), .A (n_0_0_268));
AOI21_X1 i_0_0_204 (.ZN (n_0_0_266), .A (n_0_0_275), .B1 (n_0_0_379), .B2 (n_0_0_365));
AOI21_X1 i_0_0_203 (.ZN (n_0_0_265), .A (n_0_0_266), .B1 (n_0_0_64), .B2 (n_0_0_366));
XOR2_X1 i_0_0_202 (.Z (n_0_0_264), .A (n_0_0_364), .B (n_0_0_265));
AOI22_X1 i_0_0_201 (.ZN (n_0_0_263), .A1 (n_0_0_273), .A2 (n_0_0_271), .B1 (n_0_0_269), .B2 (n_0_0_264));
OAI21_X2 i_0_0_200 (.ZN (product[14]), .A (n_0_0_263), .B1 (n_0_0_276), .B2 (n_0_0_268));
OAI22_X1 i_0_0_199 (.ZN (n_0_0_262), .A1 (n_0_0_379), .A2 (n_0_0_365), .B1 (n_0_0_64), .B2 (n_0_0_366));
AOI221_X1 i_0_0_198 (.ZN (n_0_0_261), .A (n_0_0_272), .B1 (multiplicand[6]), .B2 (n_0_0_69)
    , .C1 (n_0_0_394), .C2 (n_0_0_378));
AOI21_X1 i_0_0_197 (.ZN (n_0_0_260), .A (n_0_0_261), .B1 (n_0_0_269), .B2 (n_0_0_262));
XNOR2_X1 i_0_0_196 (.ZN (product[13]), .A (n_0_0_275), .B (n_0_0_260));
AOI22_X1 i_0_0_195 (.ZN (n_0_0_259), .A1 (n_0_0_380), .A2 (n_0_0_365), .B1 (n_0_0_54), .B2 (n_0_0_366));
OAI33_X1 i_0_0_194 (.ZN (n_0_0_258), .A1 (n_0_0_393), .A2 (multiplier[5]), .A3 (n_0_0_259)
    , .B1 (n_0_0_284), .B2 (n_0_0_283), .B3 (n_0_0_281));
XNOR2_X1 i_0_0_193 (.ZN (n_0_0_257), .A (n_0_0_291), .B (n_0_0_258));
AOI222_X1 i_0_0_192 (.ZN (n_0_0_256), .A1 (n_0_0_146), .A2 (n_0_0_273), .B1 (n_0_0_141)
    , .B2 (n_0_0_269), .C1 (n_0_0_267), .C2 (n_0_0_257));
INV_X1 i_0_0_191 (.ZN (product[12]), .A (n_0_0_256));
OAI22_X1 i_0_0_190 (.ZN (n_0_0_255), .A1 (n_0_0_44), .A2 (n_0_0_366), .B1 (n_0_0_382), .B2 (n_0_0_365));
AOI221_X1 i_0_0_189 (.ZN (n_0_0_254), .A (n_0_0_296), .B1 (n_0_0_394), .B2 (n_0_0_381)
    , .C1 (multiplicand[6]), .C2 (n_0_0_49));
AOI21_X1 i_0_0_188 (.ZN (n_0_0_253), .A (n_0_0_254), .B1 (n_0_0_361), .B2 (n_0_0_255));
XNOR2_X1 i_0_0_187 (.ZN (n_0_0_252), .A (n_0_0_301), .B (n_0_0_253));
AOI222_X2 i_0_0_186 (.ZN (n_0_0_251), .A1 (n_0_0_131), .A2 (n_0_0_286), .B1 (n_0_0_136)
    , .B2 (n_0_0_280), .C1 (n_0_0_277), .C2 (n_0_0_252));
INV_X2 i_0_0_185 (.ZN (n_0_0_250), .A (n_0_0_251));
AOI22_X1 i_0_0_184 (.ZN (n_0_0_249), .A1 (n_0_0_145), .A2 (n_0_0_273), .B1 (n_0_0_140), .B2 (n_0_0_269));
OAI21_X1 i_0_0_183 (.ZN (product[11]), .A (n_0_0_249), .B1 (n_0_0_268), .B2 (n_0_0_251));
AOI22_X1 i_0_0_182 (.ZN (n_0_0_248), .A1 (n_0_0_383), .A2 (n_0_0_365), .B1 (n_0_0_34), .B2 (n_0_0_366));
OAI33_X1 i_0_0_181 (.ZN (n_0_0_247), .A1 (n_0_0_391), .A2 (multiplier[3]), .A3 (n_0_0_248)
    , .B1 (n_0_0_306), .B2 (n_0_0_305), .B3 (n_0_0_310));
XOR2_X1 i_0_0_180 (.Z (spw__n69), .A (n_0_0_314), .B (n_0_0_247));
AOI222_X1 i_0_0_179 (.ZN (spt__n28), .A1 (n_0_0_126), .A2 (n_0_0_295), .B1 (n_0_0_121)
    , .B2 (n_0_0_361), .C1 (n_0_0_292), .C2 (n_0_0_246));
INV_X2 i_0_0_178 (.ZN (n_0_0_244), .A (n_0_0_245));
AOI22_X1 i_0_0_177 (.ZN (n_0_0_243), .A1 (n_0_0_135), .A2 (n_0_0_280), .B1 (n_0_0_130), .B2 (n_0_0_286));
OAI21_X1 i_0_0_176 (.ZN (n_0_0_242), .A (n_0_0_243), .B1 (n_0_0_278), .B2 (n_0_0_245));
AOI222_X1 i_0_0_175 (.ZN (n_0_0_241), .A1 (n_0_0_144), .A2 (n_0_0_273), .B1 (n_0_0_139)
    , .B2 (n_0_0_269), .C1 (n_0_0_267), .C2 (n_0_0_242));
INV_X1 i_0_0_174 (.ZN (product[10]), .A (n_0_0_241));
AOI22_X1 i_0_0_173 (.ZN (n_0_0_240), .A1 (n_0_0_384), .A2 (n_0_0_365), .B1 (n_0_0_24), .B2 (n_0_0_366));
OAI33_X1 i_0_0_172 (.ZN (n_0_0_239), .A1 (n_0_0_390), .A2 (multiplier[2]), .A3 (n_0_0_240)
    , .B1 (n_0_0_323), .B2 (n_0_0_322), .B3 (n_0_0_320));
XNOR2_X1 i_0_0_171 (.ZN (n_0_0_238), .A (n_0_0_327), .B (n_0_0_239));
AOI222_X2 i_0_0_170 (.ZN (n_0_0_237), .A1 (n_0_0_116), .A2 (n_0_0_309), .B1 (n_0_0_111)
    , .B2 (n_0_0_359), .C1 (n_0_0_307), .C2 (n_0_0_238));
INV_X1 i_0_0_169 (.ZN (n_0_0_236), .A (n_0_0_237));
AOI22_X1 i_0_0_168 (.ZN (n_0_0_235), .A1 (n_0_0_120), .A2 (n_0_0_361), .B1 (n_0_0_125), .B2 (n_0_0_295));
OAI21_X1 i_0_0_167 (.ZN (n_0_0_234), .A (n_0_0_235), .B1 (n_0_0_293), .B2 (n_0_0_237));
AOI222_X1 i_0_0_166 (.ZN (n_0_0_233), .A1 (n_0_0_134), .A2 (n_0_0_280), .B1 (n_0_0_129)
    , .B2 (n_0_0_286), .C1 (n_0_0_277), .C2 (n_0_0_234));
INV_X1 i_0_0_165 (.ZN (n_0_0_232), .A (n_0_0_233));
AOI22_X1 i_0_0_164 (.ZN (n_0_0_231), .A1 (n_0_0_138), .A2 (n_0_0_269), .B1 (n_0_0_143), .B2 (n_0_0_273));
OAI21_X1 i_0_0_163 (.ZN (product[9]), .A (n_0_0_231), .B1 (n_0_0_268), .B2 (n_0_0_233));
AOI22_X1 i_0_0_162 (.ZN (n_0_0_230), .A1 (n_0_0_385), .A2 (n_0_0_365), .B1 (n_0_0_14), .B2 (n_0_0_366));
OAI33_X1 i_0_0_161 (.ZN (n_0_0_229), .A1 (n_0_0_389), .A2 (multiplier[1]), .A3 (n_0_0_230)
    , .B1 (n_0_0_341), .B2 (n_0_0_340), .B3 (n_0_0_338));
XOR2_X1 i_0_0_160 (.Z (spw__n66), .A (n_0_0_342), .B (n_0_0_229));
AOI222_X1 i_0_0_159 (.ZN (n_0_0_227), .A1 (n_0_0_101), .A2 (n_0_0_357), .B1 (n_0_0_106)
    , .B2 (n_0_0_319), .C1 (n_0_0_316), .C2 (n_0_0_228));
INV_X1 i_0_0_158 (.ZN (n_0_0_226), .A (n_0_0_227));
AOI22_X1 i_0_0_157 (.ZN (n_0_0_225), .A1 (n_0_0_110), .A2 (n_0_0_359), .B1 (n_0_0_115), .B2 (n_0_0_309));
OAI21_X1 i_0_0_156 (.ZN (n_0_0_224), .A (n_0_0_225), .B1 (n_0_0_308), .B2 (n_0_0_227));
AOI222_X1 i_0_0_155 (.ZN (spw__n105), .A1 (n_0_0_119), .A2 (n_0_0_361), .B1 (n_0_0_124)
    , .B2 (n_0_0_295), .C1 (n_0_0_292), .C2 (n_0_0_224));
INV_X1 i_0_0_154 (.ZN (n_0_0_222), .A (n_0_0_223));
AOI22_X1 i_0_0_153 (.ZN (n_0_0_221), .A1 (n_0_0_133), .A2 (n_0_0_280), .B1 (n_0_0_128), .B2 (n_0_0_286));
OAI21_X1 i_0_0_152 (.ZN (n_0_0_220), .A (n_0_0_221), .B1 (n_0_0_278), .B2 (n_0_0_223));
AOI222_X1 i_0_0_151 (.ZN (n_0_0_219), .A1 (n_0_0_137), .A2 (n_0_0_269), .B1 (n_0_0_142)
    , .B2 (n_0_0_273), .C1 (n_0_0_267), .C2 (n_0_0_220));
INV_X1 i_0_0_150 (.ZN (product[8]), .A (n_0_0_219));
NAND2_X1 i_0_0_149 (.ZN (n_0_0_218), .A1 (n_0_0_353), .A2 (n_0_0_352));
XNOR2_X1 i_0_0_148 (.ZN (n_0_0_217), .A (n_0_0_386), .B (n_0_0_218));
OAI22_X1 i_0_0_147 (.ZN (n_0_0_216), .A1 (n_0_0_387), .A2 (n_0_0_365), .B1 (n_0_0_6), .B2 (n_0_0_366));
AOI221_X1 i_0_0_146 (.ZN (n_0_0_215), .A (n_0_0_348), .B1 (n_0_0_345), .B2 (n_0_0_216)
    , .C1 (n_0_0_350), .C2 (n_0_0_217));
INV_X1 i_0_0_145 (.ZN (n_0_0_214), .A (n_0_0_215));
AOI22_X1 i_0_0_144 (.ZN (n_0_0_213), .A1 (n_0_0_91), .A2 (n_0_0_334), .B1 (n_0_0_96), .B2 (n_0_0_337));
OAI21_X1 i_0_0_143 (.ZN (n_0_0_212), .A (n_0_0_213), .B1 (n_0_0_333), .B2 (n_0_0_215));
AOI222_X1 i_0_0_142 (.ZN (n_0_0_211), .A1 (n_0_0_100), .A2 (n_0_0_357), .B1 (n_0_0_105)
    , .B2 (n_0_0_319), .C1 (n_0_0_316), .C2 (n_0_0_212));
INV_X1 i_0_0_141 (.ZN (n_0_0_210), .A (n_0_0_211));
AOI22_X1 i_0_0_140 (.ZN (n_0_0_209), .A1 (n_0_0_109), .A2 (n_0_0_359), .B1 (n_0_0_114), .B2 (n_0_0_309));
OAI21_X1 i_0_0_139 (.ZN (n_0_0_208), .A (n_0_0_209), .B1 (n_0_0_308), .B2 (n_0_0_211));
AOI222_X1 i_0_0_138 (.ZN (n_0_0_207), .A1 (n_0_0_118), .A2 (n_0_0_361), .B1 (n_0_0_123)
    , .B2 (n_0_0_295), .C1 (n_0_0_292), .C2 (n_0_0_208));
INV_X1 i_0_0_137 (.ZN (n_0_0_206), .A (n_0_0_207));
AOI222_X1 i_0_0_136 (.ZN (n_0_0_205), .A1 (n_0_0_132), .A2 (n_0_0_280), .B1 (n_0_0_127)
    , .B2 (n_0_0_286), .C1 (n_0_0_277), .C2 (n_0_0_206));
INV_X1 i_0_0_135 (.ZN (n_0_0_204), .A (n_0_0_205));
NOR2_X1 i_0_0_134 (.ZN (n_0_0_203), .A1 (n_0_0_153), .A2 (n_0_0_267));
AOI21_X1 i_0_0_133 (.ZN (product[7]), .A (n_0_0_203), .B1 (n_0_0_267), .B2 (n_0_0_205));
AND2_X1 i_0_0_132 (.ZN (n_0_0_202), .A1 (multiplier[1]), .A2 (multiplier[0]));
AOI222_X2 i_0_0_131 (.ZN (n_0_0_201), .A1 (n_0_0_86), .A2 (n_0_0_350), .B1 (n_0_0_81)
    , .B2 (n_0_0_345), .C1 (n_0_0_365), .C2 (n_0_0_202));
INV_X2 i_0_0_130 (.ZN (n_0_0_200), .A (n_0_0_201));
AOI22_X1 i_0_0_129 (.ZN (n_0_0_199), .A1 (n_0_0_95), .A2 (n_0_0_337), .B1 (n_0_0_90), .B2 (n_0_0_334));
OAI21_X1 i_0_0_128 (.ZN (n_0_0_198), .A (n_0_0_199), .B1 (n_0_0_333), .B2 (n_0_0_201));
AOI222_X1 i_0_0_127 (.ZN (n_0_0_197), .A1 (n_0_0_99), .A2 (n_0_0_357), .B1 (n_0_0_104)
    , .B2 (n_0_0_319), .C1 (n_0_0_316), .C2 (n_0_0_198));
INV_X1 i_0_0_126 (.ZN (n_0_0_196), .A (n_0_0_197));
AOI22_X1 i_0_0_125 (.ZN (n_0_0_195), .A1 (n_0_0_108), .A2 (n_0_0_359), .B1 (n_0_0_113), .B2 (n_0_0_309));
OAI21_X1 i_0_0_124 (.ZN (n_0_0_194), .A (n_0_0_195), .B1 (n_0_0_308), .B2 (n_0_0_197));
AOI222_X1 i_0_0_123 (.ZN (n_0_0_193), .A1 (n_0_0_117), .A2 (n_0_0_361), .B1 (n_0_0_122)
    , .B2 (n_0_0_295), .C1 (n_0_0_292), .C2 (n_0_0_194));
INV_X1 i_0_0_122 (.ZN (n_0_0_192), .A (n_0_0_193));
NOR2_X1 i_0_0_121 (.ZN (n_0_0_191), .A1 (n_0_0_152), .A2 (n_0_0_277));
AOI21_X1 i_0_0_120 (.ZN (product[6]), .A (n_0_0_191), .B1 (n_0_0_277), .B2 (n_0_0_193));
AOI21_X2 i_0_0_119 (.ZN (spt__n36), .A (n_0_0_369), .B1 (multiplicand[5]), .B2 (n_0_0_370));
AOI222_X2 i_0_0_118 (.ZN (n_0_0_189), .A1 (n_0_0_80), .A2 (n_0_0_345), .B1 (n_0_0_85)
    , .B2 (n_0_0_350), .C1 (n_0_0_202), .C2 (n_0_0_190));
INV_X2 i_0_0_117 (.ZN (n_0_0_188), .A (n_0_0_189));
AOI22_X1 i_0_0_116 (.ZN (n_0_0_187), .A1 (n_0_0_94), .A2 (n_0_0_337), .B1 (n_0_0_89), .B2 (n_0_0_334));
OAI21_X1 i_0_0_115 (.ZN (n_0_0_186), .A (n_0_0_187), .B1 (n_0_0_333), .B2 (n_0_0_189));
AOI222_X1 i_0_0_114 (.ZN (n_0_0_185), .A1 (n_0_0_98), .A2 (n_0_0_357), .B1 (n_0_0_103)
    , .B2 (n_0_0_319), .C1 (n_0_0_316), .C2 (n_0_0_186));
INV_X1 i_0_0_113 (.ZN (n_0_0_184), .A (n_0_0_185));
AOI222_X1 i_0_0_112 (.ZN (n_0_0_183), .A1 (n_0_0_107), .A2 (n_0_0_359), .B1 (n_0_0_112)
    , .B2 (n_0_0_309), .C1 (n_0_0_307), .C2 (n_0_0_184));
INV_X1 i_0_0_111 (.ZN (n_0_0_182), .A (n_0_0_183));
NOR2_X1 i_0_0_110 (.ZN (n_0_0_181), .A1 (n_0_0_151), .A2 (n_0_0_292));
AOI21_X1 i_0_0_109 (.ZN (product[5]), .A (n_0_0_181), .B1 (n_0_0_292), .B2 (n_0_0_183));
AOI21_X2 i_0_0_108 (.ZN (spt__n41), .A (n_0_0_371), .B1 (multiplicand[4]), .B2 (n_0_0_372));
AOI222_X2 i_0_0_107 (.ZN (n_0_0_179), .A1 (n_0_0_79), .A2 (n_0_0_345), .B1 (n_0_0_84)
    , .B2 (n_0_0_350), .C1 (n_0_0_202), .C2 (n_0_0_180));
INV_X2 i_0_0_106 (.ZN (n_0_0_178), .A (n_0_0_179));
AOI22_X1 i_0_0_105 (.ZN (n_0_0_177), .A1 (n_0_0_88), .A2 (n_0_0_334), .B1 (n_0_0_93), .B2 (n_0_0_337));
OAI21_X1 i_0_0_104 (.ZN (n_0_0_176), .A (n_0_0_177), .B1 (n_0_0_333), .B2 (n_0_0_179));
AOI222_X1 i_0_0_103 (.ZN (n_0_0_175), .A1 (n_0_0_97), .A2 (n_0_0_357), .B1 (n_0_0_102)
    , .B2 (n_0_0_319), .C1 (n_0_0_316), .C2 (n_0_0_176));
INV_X1 i_0_0_102 (.ZN (n_0_0_174), .A (n_0_0_175));
NOR2_X1 i_0_0_101 (.ZN (n_0_0_173), .A1 (n_0_0_150), .A2 (n_0_0_307));
AOI21_X1 i_0_0_100 (.ZN (product[4]), .A (n_0_0_173), .B1 (n_0_0_307), .B2 (n_0_0_175));
AOI21_X1 i_0_0_99 (.ZN (spt__n31), .A (n_0_0_373), .B1 (multiplicand[3]), .B2 (n_0_0_374));
AOI222_X2 i_0_0_98 (.ZN (n_0_0_171), .A1 (n_0_0_83), .A2 (n_0_0_350), .B1 (n_0_0_78)
    , .B2 (n_0_0_345), .C1 (n_0_0_202), .C2 (spw__n692));
INV_X2 i_0_0_97 (.ZN (n_0_0_170), .A (n_0_0_171));
AOI22_X1 i_0_0_96 (.ZN (n_0_0_169), .A1 (n_0_0_92), .A2 (n_0_0_337), .B1 (n_0_0_87), .B2 (n_0_0_334));
OAI21_X1 i_0_0_95 (.ZN (n_0_0_168), .A (n_0_0_169), .B1 (n_0_0_333), .B2 (n_0_0_171));
AOI22_X1 i_0_0_94 (.ZN (n_0_0_167), .A1 (n_0_0_149), .A2 (n_0_0_317), .B1 (n_0_0_316), .B2 (n_0_0_168));
INV_X1 i_0_0_93 (.ZN (product[3]), .A (n_0_0_167));
AOI21_X4 i_0_0_92 (.ZN (n_0_0_166), .A (n_0_0_375), .B1 (multiplicand[2]), .B2 (n_0_0_376));
AOI222_X1 i_0_0_91 (.ZN (n_0_0_165), .A1 (n_0_0_82), .A2 (n_0_0_350), .B1 (n_0_0_77)
    , .B2 (n_0_0_345), .C1 (n_0_0_202), .C2 (spw__n582));
INV_X1 i_0_0_90 (.ZN (n_0_0_164), .A (n_0_0_165));
NAND2_X1 i_0_0_89 (.ZN (n_0_0_163), .A1 (n_0_0_148), .A2 (n_0_0_333));
OAI21_X1 i_0_0_88 (.ZN (product[2]), .A (n_0_0_163), .B1 (n_0_0_333), .B2 (n_0_0_165));
OAI21_X1 i_0_0_87 (.ZN (n_0_0_162), .A (n_0_0_147), .B1 (n_0_0_350), .B2 (n_0_0_345));
AOI21_X2 i_0_0_86 (.ZN (n_0_0_161), .A (n_0_0_377), .B1 (multiplicand[1]), .B2 (multiplicand[0]));
NAND2_X4 i_0_0_85 (.ZN (n_0_0_160), .A1 (multiplier[0]), .A2 (spc__n4));
INV_X4 i_0_0_84 (.ZN (n_0_0_159), .A (n_0_0_160));
OAI21_X1 i_0_0_83 (.ZN (product[1]), .A (n_0_0_162), .B1 (n_0_0_388), .B2 (spw__n662));
AND2_X1 i_0_0_82 (.ZN (product[0]), .A1 (spw__n165), .A2 (multiplier[0]));
AND2_X1 i_0_0_81 (.ZN (n_0_0_158), .A1 (multiplier[0]), .A2 (n_0_0_166));
AND2_X4 i_0_0_80 (.ZN (n_0_0_157), .A1 (multiplier[0]), .A2 (n_0_0_172));
AND2_X4 i_0_0_79 (.ZN (n_0_0_156), .A1 (multiplier[0]), .A2 (n_0_0_180));
AND2_X4 i_0_0_78 (.ZN (n_0_0_155), .A1 (multiplier[0]), .A2 (n_0_0_190));
AND2_X1 i_0_0_77 (.ZN (n_0_0_154), .A1 (multiplier[0]), .A2 (n_0_0_365));
HA_X1 i_0_0_76 (.CO (n_0_0_76), .S (n_0_0_153), .A (spw__n162), .B (n_0_0_204));
HA_X1 i_0_0_75 (.CO (n_0_0_75), .S (n_0_0_152), .A (spw__n165), .B (n_0_0_192));
HA_X1 i_0_0_74 (.CO (n_0_0_74), .S (n_0_0_151), .A (spw__n165), .B (n_0_0_182));
HA_X1 i_0_0_73 (.CO (n_0_0_73), .S (n_0_0_150), .A (spw__n164), .B (n_0_0_174));
HA_X1 i_0_0_72 (.CO (n_0_0_72), .S (n_0_0_149), .A (spw__n164), .B (n_0_0_168));
HA_X1 i_0_0_71 (.CO (n_0_0_71), .S (n_0_0_148), .A (spw__n166), .B (n_0_0_164));
HA_X1 i_0_0_70 (.CO (n_0_0_70), .S (n_0_0_147), .A (spw__n163), .B (n_0_0_159));
FA_X1 i_0_0_69 (.CO (n_0_0_69), .S (n_0_0_146), .A (multiplicand[5]), .B (n_0_0_257), .CI (n_0_0_68));
FA_X1 i_0_0_68 (.CO (n_0_0_68), .S (n_0_0_145), .A (multiplicand[4]), .B (n_0_0_250), .CI (n_0_0_67));
FA_X1 i_0_0_67 (.CO (n_0_0_67), .S (n_0_0_144), .A (multiplicand[3]), .B (n_0_0_242), .CI (n_0_0_66));
FA_X1 i_0_0_66 (.CO (n_0_0_66), .S (n_0_0_143), .A (multiplicand[2]), .B (n_0_0_232), .CI (n_0_0_65));
FA_X1 i_0_0_65 (.CO (n_0_0_65), .S (n_0_0_142), .A (multiplicand[1]), .B (n_0_0_220), .CI (n_0_0_76));
FA_X1 i_0_0_64 (.CO (n_0_0_64), .S (n_0_0_141), .A (n_0_0_190), .B (n_0_0_257), .CI (n_0_0_63));
FA_X1 i_0_0_63 (.CO (n_0_0_63), .S (n_0_0_140), .A (n_0_0_180), .B (n_0_0_250), .CI (n_0_0_62));
FA_X1 i_0_0_62 (.CO (n_0_0_62), .S (n_0_0_139), .A (spw__n683), .B (n_0_0_242), .CI (n_0_0_61));
FA_X1 i_0_0_61 (.CO (n_0_0_61), .S (n_0_0_138), .A (spw__n584), .B (n_0_0_232), .CI (n_0_0_60));
FA_X1 i_0_0_60 (.CO (n_0_0_60), .S (n_0_0_137), .A (spc__n9), .B (n_0_0_220), .CI (n_0_0_76));
FA_X1 i_0_0_59 (.CO (n_0_0_59), .S (n_0_0_136), .A (multiplicand[5]), .B (n_0_0_252), .CI (n_0_0_58));
FA_X1 i_0_0_58 (.CO (n_0_0_58), .S (n_0_0_135), .A (multiplicand[4]), .B (n_0_0_244), .CI (n_0_0_57));
FA_X1 i_0_0_57 (.CO (n_0_0_57), .S (n_0_0_134), .A (multiplicand[3]), .B (n_0_0_234), .CI (n_0_0_56));
FA_X1 i_0_0_56 (.CO (n_0_0_56), .S (n_0_0_133), .A (multiplicand[2]), .B (n_0_0_222), .CI (n_0_0_55));
FA_X1 i_0_0_55 (.CO (n_0_0_55), .S (n_0_0_132), .A (multiplicand[1]), .B (n_0_0_206), .CI (n_0_0_75));
FA_X1 i_0_0_54 (.CO (n_0_0_54), .S (n_0_0_131), .A (n_0_0_190), .B (n_0_0_252), .CI (n_0_0_53));
FA_X1 i_0_0_53 (.CO (n_0_0_53), .S (n_0_0_130), .A (n_0_0_180), .B (n_0_0_244), .CI (n_0_0_52));
FA_X1 i_0_0_52 (.CO (n_0_0_52), .S (n_0_0_129), .A (spw__n684), .B (n_0_0_234), .CI (n_0_0_51));
FA_X1 i_0_0_51 (.CO (n_0_0_51), .S (n_0_0_128), .A (spw__n577), .B (n_0_0_222), .CI (n_0_0_50));
FA_X1 i_0_0_50 (.CO (n_0_0_50), .S (n_0_0_127), .A (spc__n8), .B (n_0_0_206), .CI (n_0_0_75));
FA_X1 i_0_0_49 (.CO (n_0_0_49), .S (n_0_0_126), .A (multiplicand[5]), .B (n_0_0_246), .CI (n_0_0_48));
FA_X1 i_0_0_48 (.CO (n_0_0_48), .S (n_0_0_125), .A (multiplicand[4]), .B (n_0_0_236), .CI (n_0_0_47));
FA_X1 i_0_0_47 (.CO (n_0_0_47), .S (n_0_0_124), .A (multiplicand[3]), .B (n_0_0_224), .CI (n_0_0_46));
FA_X1 i_0_0_46 (.CO (n_0_0_46), .S (n_0_0_123), .A (multiplicand[2]), .B (n_0_0_208), .CI (n_0_0_45));
FA_X1 i_0_0_45 (.CO (n_0_0_45), .S (n_0_0_122), .A (multiplicand[1]), .B (n_0_0_194), .CI (n_0_0_74));
FA_X1 i_0_0_44 (.CO (n_0_0_44), .S (n_0_0_121), .A (n_0_0_190), .B (n_0_0_246), .CI (n_0_0_43));
FA_X1 i_0_0_43 (.CO (n_0_0_43), .S (n_0_0_120), .A (n_0_0_180), .B (n_0_0_236), .CI (n_0_0_42));
FA_X1 i_0_0_42 (.CO (n_0_0_42), .S (n_0_0_119), .A (spw__n686), .B (n_0_0_224), .CI (n_0_0_41));
FA_X1 i_0_0_41 (.CO (n_0_0_41), .S (n_0_0_118), .A (spw__n578), .B (n_0_0_208), .CI (n_0_0_40));
FA_X1 i_0_0_40 (.CO (n_0_0_40), .S (n_0_0_117), .A (spc__n7), .B (n_0_0_194), .CI (n_0_0_74));
FA_X1 i_0_0_39 (.CO (n_0_0_39), .S (n_0_0_116), .A (multiplicand[5]), .B (n_0_0_238), .CI (n_0_0_38));
FA_X1 i_0_0_38 (.CO (n_0_0_38), .S (n_0_0_115), .A (multiplicand[4]), .B (n_0_0_226), .CI (n_0_0_37));
FA_X1 i_0_0_37 (.CO (n_0_0_37), .S (n_0_0_114), .A (multiplicand[3]), .B (n_0_0_210), .CI (n_0_0_36));
FA_X1 i_0_0_36 (.CO (n_0_0_36), .S (n_0_0_113), .A (multiplicand[2]), .B (n_0_0_196), .CI (n_0_0_35));
FA_X1 i_0_0_35 (.CO (n_0_0_35), .S (n_0_0_112), .A (multiplicand[1]), .B (n_0_0_184), .CI (n_0_0_73));
FA_X1 i_0_0_34 (.CO (n_0_0_34), .S (n_0_0_111), .A (n_0_0_190), .B (n_0_0_238), .CI (n_0_0_33));
FA_X1 i_0_0_33 (.CO (n_0_0_33), .S (n_0_0_110), .A (n_0_0_180), .B (n_0_0_226), .CI (n_0_0_32));
FA_X1 i_0_0_32 (.CO (n_0_0_32), .S (n_0_0_109), .A (spw__n687), .B (n_0_0_210), .CI (n_0_0_31));
FA_X1 i_0_0_31 (.CO (n_0_0_31), .S (n_0_0_108), .A (spw__n579), .B (n_0_0_196), .CI (n_0_0_30));
FA_X1 i_0_0_30 (.CO (n_0_0_30), .S (n_0_0_107), .A (spc__n2), .B (n_0_0_184), .CI (n_0_0_73));
FA_X1 i_0_0_29 (.CO (n_0_0_29), .S (n_0_0_106), .A (multiplicand[5]), .B (n_0_0_228), .CI (n_0_0_28));
FA_X1 i_0_0_28 (.CO (n_0_0_28), .S (n_0_0_105), .A (multiplicand[4]), .B (n_0_0_212), .CI (n_0_0_27));
FA_X1 i_0_0_27 (.CO (n_0_0_27), .S (n_0_0_104), .A (multiplicand[3]), .B (n_0_0_198), .CI (n_0_0_26));
FA_X1 i_0_0_26 (.CO (n_0_0_26), .S (n_0_0_103), .A (multiplicand[2]), .B (n_0_0_186), .CI (n_0_0_25));
FA_X1 i_0_0_25 (.CO (n_0_0_25), .S (n_0_0_102), .A (multiplicand[1]), .B (n_0_0_176), .CI (n_0_0_72));
FA_X1 i_0_0_24 (.CO (n_0_0_24), .S (n_0_0_101), .A (n_0_0_190), .B (n_0_0_228), .CI (n_0_0_23));
FA_X1 i_0_0_23 (.CO (n_0_0_23), .S (n_0_0_100), .A (n_0_0_180), .B (n_0_0_212), .CI (n_0_0_22));
FA_X1 i_0_0_22 (.CO (n_0_0_22), .S (n_0_0_99), .A (spw__n688), .B (n_0_0_198), .CI (n_0_0_21));
FA_X1 i_0_0_21 (.CO (n_0_0_21), .S (n_0_0_98), .A (spw__n580), .B (n_0_0_186), .CI (n_0_0_20));
FA_X1 i_0_0_20 (.CO (n_0_0_20), .S (n_0_0_97), .A (spc__n3), .B (n_0_0_176), .CI (n_0_0_72));
FA_X1 i_0_0_19 (.CO (n_0_0_19), .S (n_0_0_96), .A (multiplicand[5]), .B (n_0_0_214), .CI (n_0_0_18));
FA_X1 i_0_0_18 (.CO (n_0_0_18), .S (n_0_0_95), .A (multiplicand[4]), .B (n_0_0_200), .CI (n_0_0_17));
FA_X1 i_0_0_17 (.CO (n_0_0_17), .S (n_0_0_94), .A (multiplicand[3]), .B (n_0_0_188), .CI (n_0_0_16));
FA_X1 i_0_0_16 (.CO (n_0_0_16), .S (n_0_0_93), .A (multiplicand[2]), .B (n_0_0_178), .CI (n_0_0_15));
FA_X1 i_0_0_15 (.CO (n_0_0_15), .S (n_0_0_92), .A (multiplicand[1]), .B (n_0_0_170), .CI (n_0_0_71));
FA_X1 i_0_0_14 (.CO (n_0_0_14), .S (n_0_0_91), .A (n_0_0_190), .B (n_0_0_214), .CI (n_0_0_13));
FA_X1 i_0_0_13 (.CO (n_0_0_13), .S (n_0_0_90), .A (n_0_0_180), .B (n_0_0_200), .CI (n_0_0_12));
FA_X1 i_0_0_12 (.CO (n_0_0_12), .S (n_0_0_89), .A (spw__n691), .B (n_0_0_188), .CI (n_0_0_11));
FA_X1 i_0_0_11 (.CO (n_0_0_11), .S (n_0_0_88), .A (spw__n581), .B (n_0_0_178), .CI (n_0_0_10));
FA_X1 i_0_0_10 (.CO (n_0_0_10), .S (n_0_0_87), .A (spc__n6), .B (n_0_0_170), .CI (n_0_0_71));
FA_X1 i_0_0_9 (.CO (n_0_0_9), .S (n_0_0_86), .A (multiplicand[5]), .B (n_0_0_154), .CI (n_0_0_8));
FA_X1 i_0_0_8 (.CO (n_0_0_8), .S (n_0_0_85), .A (multiplicand[4]), .B (n_0_0_155), .CI (n_0_0_7));
FA_X1 i_0_0_7 (.CO (n_0_0_7), .S (n_0_0_84), .A (multiplicand[3]), .B (n_0_0_156), .CI (n_0_0_1));
FA_X1 i_0_0_6 (.CO (n_0_0_1), .S (n_0_0_83), .A (multiplicand[2]), .B (n_0_0_157), .CI (n_0_0_0));
FA_X1 i_0_0_5 (.CO (n_0_0_0), .S (n_0_0_82), .A (multiplicand[1]), .B (n_0_0_158), .CI (n_0_0_70));
FA_X1 i_0_0_4 (.CO (n_0_0_6), .S (n_0_0_81), .A (n_0_0_190), .B (n_0_0_154), .CI (n_0_0_5));
FA_X1 i_0_0_3 (.CO (n_0_0_5), .S (n_0_0_80), .A (n_0_0_180), .B (n_0_0_155), .CI (n_0_0_4));
FA_X1 i_0_0_2 (.CO (n_0_0_4), .S (n_0_0_79), .A (spw__n689), .B (n_0_0_156), .CI (n_0_0_3));
FA_X1 i_0_0_1 (.CO (n_0_0_3), .S (n_0_0_78), .A (spw__n583), .B (n_0_0_157), .CI (n_0_0_2));
FA_X1 i_0_0_0 (.CO (n_0_0_2), .S (n_0_0_77), .A (spc__n5), .B (n_0_0_158), .CI (n_0_0_70));
BUF_X4 spc__L1_c1 (.Z (spc__n1), .A (n_0_0_161));
BUF_X1 spc__L2_c2 (.Z (spc__n2), .A (spc__n1));
BUF_X1 spc__L2_c3 (.Z (spc__n3), .A (spc__n1));
BUF_X4 spc__L2_c4 (.Z (spc__n4), .A (spc__n1));
BUF_X2 spc__L2_c5 (.Z (spc__n5), .A (spc__n1));
BUF_X1 spc__L2_c6 (.Z (spc__n6), .A (spc__n1));
BUF_X1 spc__L2_c7 (.Z (spc__n7), .A (spc__n1));
BUF_X2 spc__L2_c8 (.Z (spc__n8), .A (spc__n1));
BUF_X1 spc__L2_c9 (.Z (spc__n9), .A (spc__n1));
BUF_X1 spt__c28 (.Z (n_0_0_245), .A (spt__n28));
BUF_X4 spt__c31 (.Z (n_0_0_172), .A (spt__n31));
BUF_X4 spt__c36 (.Z (n_0_0_190), .A (spt__n36));
BUF_X4 spt__c41 (.Z (n_0_0_180), .A (spt__n41));
BUF_X4 spw__c64 (.Z (n_0_0_228), .A (spw__n66));
BUF_X2 spw__c67 (.Z (n_0_0_246), .A (spw__n69));
CLKBUF_X2 spw__c103 (.Z (n_0_0_223), .A (spw__n105));
BUF_X1 spw__L1_c160 (.Z (spw__n162), .A (multiplicand[0]));
BUF_X1 spw__L1_c161 (.Z (spw__n163), .A (multiplicand[0]));
BUF_X1 spw__L2_c162 (.Z (spw__n164), .A (spw__n163));
BUF_X2 spw__L3_c163 (.Z (spw__n165), .A (spw__n164));
BUF_X1 spw__L2_c164 (.Z (spw__n166), .A (spw__n163));
INV_X1 spw__L1_c568 (.ZN (spw__n572), .A (n_0_0_166));
BUF_X1 spw__L2_c569 (.Z (spw__n573), .A (spw__n572));
BUF_X1 spw__L3_c570 (.Z (spw__n574), .A (spw__n573));
BUF_X1 spw__L4_c571 (.Z (spw__n575), .A (spw__n574));
BUF_X1 spw__L5_c572 (.Z (spw__n576), .A (spw__n575));
INV_X1 spw__L6_c573 (.ZN (spw__n577), .A (spw__n576));
INV_X1 spw__L5_c574 (.ZN (spw__n578), .A (spw__n575));
INV_X1 spw__L4_c575 (.ZN (spw__n579), .A (spw__n574));
INV_X1 spw__L3_c576 (.ZN (spw__n580), .A (spw__n573));
INV_X2 spw__L2_c577 (.ZN (spw__n581), .A (spw__n572));
BUF_X1 spw__L1_c578 (.Z (spw__n582), .A (n_0_0_166));
BUF_X2 spw__L1_c579 (.Z (spw__n583), .A (n_0_0_166));
BUF_X1 spw__L1_c580 (.Z (spw__n584), .A (n_0_0_166));
CLKBUF_X1 spw__L1_c658 (.Z (spw__n662), .A (n_0_0_160));
INV_X1 spw__L1_c678 (.ZN (spw__n682), .A (n_0_0_172));
INV_X1 spw__L2_c679 (.ZN (spw__n683), .A (spw__n682));
INV_X1 spw__L2_c680 (.ZN (spw__n684), .A (spw__n682));
INV_X1 spw__L1_c681 (.ZN (spw__n685), .A (n_0_0_172));
INV_X1 spw__L2_c682 (.ZN (spw__n686), .A (spw__n685));
INV_X2 spw__L2_c683 (.ZN (spw__n687), .A (spw__n685));
BUF_X1 spw__L1_c684 (.Z (spw__n688), .A (n_0_0_172));
BUF_X2 spw__L1_c685 (.Z (spw__n689), .A (n_0_0_172));
INV_X1 spw__L1_c686 (.ZN (spw__n690), .A (n_0_0_172));
INV_X1 spw__L2_c687 (.ZN (spw__n691), .A (spw__n690));
INV_X1 spw__L2_c688 (.ZN (spw__n692), .A (spw__n690));

endmodule //Booth_Multiplier


