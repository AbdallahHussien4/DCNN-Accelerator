/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Wed May 26 17:39:58 2021
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 3487642794 */

module RAM(enable, clk, address, write, \output_data[0][0] , \output_data[0][1] , 
      \output_data[0][2] , \output_data[0][3] , \output_data[0][4] , 
      \output_data[1][0] , \output_data[1][1] , \output_data[1][2] , 
      \output_data[1][3] , \output_data[1][4] , \output_data[2][0] , 
      \output_data[2][1] , \output_data[2][2] , \output_data[2][3] , 
      \output_data[2][4] , \output_data[3][0] , \output_data[3][1] , 
      \output_data[3][2] , \output_data[3][3] , \output_data[3][4] , 
      \output_data[4][0] , \output_data[4][1] , \output_data[4][2] , 
      \output_data[4][3] , \output_data[4][4] , offset, input_data, finish);
   input enable;
   input clk;
   input [15:0]address;
   input write;
   output [15:0]\output_data[0][0] ;
   output [15:0]\output_data[0][1] ;
   output [15:0]\output_data[0][2] ;
   output [15:0]\output_data[0][3] ;
   output [15:0]\output_data[0][4] ;
   output [15:0]\output_data[1][0] ;
   output [15:0]\output_data[1][1] ;
   output [15:0]\output_data[1][2] ;
   output [15:0]\output_data[1][3] ;
   output [15:0]\output_data[1][4] ;
   output [15:0]\output_data[2][0] ;
   output [15:0]\output_data[2][1] ;
   output [15:0]\output_data[2][2] ;
   output [15:0]\output_data[2][3] ;
   output [15:0]\output_data[2][4] ;
   output [15:0]\output_data[3][0] ;
   output [15:0]\output_data[3][1] ;
   output [15:0]\output_data[3][2] ;
   output [15:0]\output_data[3][3] ;
   output [15:0]\output_data[3][4] ;
   output [15:0]\output_data[4][0] ;
   output [15:0]\output_data[4][1] ;
   output [15:0]\output_data[4][2] ;
   output [15:0]\output_data[4][3] ;
   output [15:0]\output_data[4][4] ;
   input [15:0]offset;
   input [15:0]input_data;
   output finish;

   wire n_28_0;

   DFF_X1 finish_flag_reg__0 (.D(1'b0), .CK(n_28_0), .Q(1'b0), .QN());
   INV_X1 i_28_0_0 (.A(clk), .ZN(n_28_0));
endmodule

module DMA(start, reset, finish_read, clk, address, offset, 
      read_write_filter_bias, filter_number, \CNN_output_data[0][0] , 
      \CNN_output_data[0][1] , \CNN_output_data[0][2] , \CNN_output_data[0][3] , 
      \CNN_output_data[0][4] , \CNN_output_data[1][0] , \CNN_output_data[1][1] , 
      \CNN_output_data[1][2] , \CNN_output_data[1][3] , \CNN_output_data[1][4] , 
      \CNN_output_data[2][0] , \CNN_output_data[2][1] , \CNN_output_data[2][2] , 
      \CNN_output_data[2][3] , \CNN_output_data[2][4] , \CNN_output_data[3][0] , 
      \CNN_output_data[3][1] , \CNN_output_data[3][2] , \CNN_output_data[3][3] , 
      \CNN_output_data[3][4] , \CNN_output_data[4][0] , \CNN_output_data[4][1] , 
      \CNN_output_data[4][2] , \CNN_output_data[4][3] , \CNN_output_data[4][4] , 
      CNN_input_data, RAM_address, RAM_offset, RAM_write, RAM_output_data, 
      \RAM_input_data[0][0] , \RAM_input_data[0][1] , \RAM_input_data[0][2] , 
      \RAM_input_data[0][3] , \RAM_input_data[0][4] , \RAM_input_data[1][0] , 
      \RAM_input_data[1][1] , \RAM_input_data[1][2] , \RAM_input_data[1][3] , 
      \RAM_input_data[1][4] , \RAM_input_data[2][0] , \RAM_input_data[2][1] , 
      \RAM_input_data[2][2] , \RAM_input_data[2][3] , \RAM_input_data[2][4] , 
      \RAM_input_data[3][0] , \RAM_input_data[3][1] , \RAM_input_data[3][2] , 
      \RAM_input_data[3][3] , \RAM_input_data[3][4] , \RAM_input_data[4][0] , 
      \RAM_input_data[4][1] , \RAM_input_data[4][2] , \RAM_input_data[4][3] , 
      \RAM_input_data[4][4] , RAM_finish, RAM_enable, FB_write, 
      \FB_filter[0][0] , \FB_filter[0][1] , \FB_filter[0][2] , \FB_filter[0][3] , 
      \FB_filter[0][4] , \FB_filter[1][0] , \FB_filter[1][1] , \FB_filter[1][2] , 
      \FB_filter[1][3] , \FB_filter[1][4] , \FB_filter[2][0] , \FB_filter[2][1] , 
      \FB_filter[2][2] , \FB_filter[2][3] , \FB_filter[2][4] , \FB_filter[3][0] , 
      \FB_filter[3][1] , \FB_filter[3][2] , \FB_filter[3][3] , \FB_filter[3][4] , 
      \FB_filter[4][0] , \FB_filter[4][1] , \FB_filter[4][2] , \FB_filter[4][3] , 
      \FB_filter[4][4] , FB_index_filter, \FB_bias[0] , \FB_bias[1] , 
      \FB_bias[2] , \FB_bias[3] , \FB_bias[4] , \FB_bias[5] , \FB_bias[6] , 
      \FB_bias[7] , \FB_bias[8] , \FB_bias[9] , \FB_bias[10] , \FB_bias[11] , 
      \FB_bias[12] , \FB_bias[13] , \FB_bias[14] , \FB_bias[15] , \FB_bias[16] , 
      \FB_bias[17] , \FB_bias[18] , \FB_bias[19] , \FB_bias[20] , \FB_bias[21] , 
      \FB_bias[22] , \FB_bias[23] , \FB_bias[24] , \FB_bias[25] , \FB_bias[26] , 
      \FB_bias[27] , \FB_bias[28] , \FB_bias[29] , \FB_bias[30] , \FB_bias[31] , 
      \FB_bias[32] , \FB_bias[33] , \FB_bias[34] , \FB_bias[35] , \FB_bias[36] , 
      \FB_bias[37] , \FB_bias[38] , \FB_bias[39] , \FB_bias[40] , \FB_bias[41] , 
      \FB_bias[42] , \FB_bias[43] , \FB_bias[44] , \FB_bias[45] , \FB_bias[46] , 
      \FB_bias[47] , \FB_bias[48] , \FB_bias[49] , \FB_bias[50] , \FB_bias[51] , 
      \FB_bias[52] , \FB_bias[53] , \FB_bias[54] , \FB_bias[55] , \FB_bias[56] , 
      \FB_bias[57] , \FB_bias[58] , \FB_bias[59] , \FB_bias[60] , \FB_bias[61] , 
      \FB_bias[62] , \FB_bias[63] , \FB_bias[64] , \FB_bias[65] , \FB_bias[66] , 
      \FB_bias[67] , \FB_bias[68] , \FB_bias[69] , \FB_bias[70] , \FB_bias[71] , 
      \FB_bias[72] , \FB_bias[73] , \FB_bias[74] , \FB_bias[75] , \FB_bias[76] , 
      \FB_bias[77] , \FB_bias[78] , \FB_bias[79] , \FB_bias[80] , \FB_bias[81] , 
      \FB_bias[82] , \FB_bias[83] , \FB_bias[84] , \FB_bias[85] , \FB_bias[86] , 
      \FB_bias[87] , \FB_bias[88] , \FB_bias[89] , \FB_bias[90] , \FB_bias[91] , 
      \FB_bias[92] , \FB_bias[93] , \FB_bias[94] , \FB_bias[95] , \FB_bias[96] , 
      \FB_bias[97] , \FB_bias[98] , \FB_bias[99] , \FB_bias[100] , 
      \FB_bias[101] , \FB_bias[102] , \FB_bias[103] , \FB_bias[104] , 
      \FB_bias[105] , \FB_bias[106] , \FB_bias[107] , \FB_bias[108] , 
      \FB_bias[109] , \FB_bias[110] , \FB_bias[111] , \FB_bias[112] , 
      \FB_bias[113] , \FB_bias[114] , \FB_bias[115] , \FB_bias[116] , 
      \FB_bias[117] , \FB_bias[118] , \FB_bias[119] , FB_bias_or_filter, 
      FB_finish);
   input start;
   input reset;
   output finish_read;
   input clk;
   input [15:0]address;
   input [15:0]offset;
   input [1:0]read_write_filter_bias;
   input [15:0]filter_number;
   output [15:0]\CNN_output_data[0][0] ;
   output [15:0]\CNN_output_data[0][1] ;
   output [15:0]\CNN_output_data[0][2] ;
   output [15:0]\CNN_output_data[0][3] ;
   output [15:0]\CNN_output_data[0][4] ;
   output [15:0]\CNN_output_data[1][0] ;
   output [15:0]\CNN_output_data[1][1] ;
   output [15:0]\CNN_output_data[1][2] ;
   output [15:0]\CNN_output_data[1][3] ;
   output [15:0]\CNN_output_data[1][4] ;
   output [15:0]\CNN_output_data[2][0] ;
   output [15:0]\CNN_output_data[2][1] ;
   output [15:0]\CNN_output_data[2][2] ;
   output [15:0]\CNN_output_data[2][3] ;
   output [15:0]\CNN_output_data[2][4] ;
   output [15:0]\CNN_output_data[3][0] ;
   output [15:0]\CNN_output_data[3][1] ;
   output [15:0]\CNN_output_data[3][2] ;
   output [15:0]\CNN_output_data[3][3] ;
   output [15:0]\CNN_output_data[3][4] ;
   output [15:0]\CNN_output_data[4][0] ;
   output [15:0]\CNN_output_data[4][1] ;
   output [15:0]\CNN_output_data[4][2] ;
   output [15:0]\CNN_output_data[4][3] ;
   output [15:0]\CNN_output_data[4][4] ;
   input [15:0]CNN_input_data;
   output [15:0]RAM_address;
   output [15:0]RAM_offset;
   output RAM_write;
   output [15:0]RAM_output_data;
   input [15:0]\RAM_input_data[0][0] ;
   input [15:0]\RAM_input_data[0][1] ;
   input [15:0]\RAM_input_data[0][2] ;
   input [15:0]\RAM_input_data[0][3] ;
   input [15:0]\RAM_input_data[0][4] ;
   input [15:0]\RAM_input_data[1][0] ;
   input [15:0]\RAM_input_data[1][1] ;
   input [15:0]\RAM_input_data[1][2] ;
   input [15:0]\RAM_input_data[1][3] ;
   input [15:0]\RAM_input_data[1][4] ;
   input [15:0]\RAM_input_data[2][0] ;
   input [15:0]\RAM_input_data[2][1] ;
   input [15:0]\RAM_input_data[2][2] ;
   input [15:0]\RAM_input_data[2][3] ;
   input [15:0]\RAM_input_data[2][4] ;
   input [15:0]\RAM_input_data[3][0] ;
   input [15:0]\RAM_input_data[3][1] ;
   input [15:0]\RAM_input_data[3][2] ;
   input [15:0]\RAM_input_data[3][3] ;
   input [15:0]\RAM_input_data[3][4] ;
   input [15:0]\RAM_input_data[4][0] ;
   input [15:0]\RAM_input_data[4][1] ;
   input [15:0]\RAM_input_data[4][2] ;
   input [15:0]\RAM_input_data[4][3] ;
   input [15:0]\RAM_input_data[4][4] ;
   input RAM_finish;
   output RAM_enable;
   output FB_write;
   output [15:0]\FB_filter[0][0] ;
   output [15:0]\FB_filter[0][1] ;
   output [15:0]\FB_filter[0][2] ;
   output [15:0]\FB_filter[0][3] ;
   output [15:0]\FB_filter[0][4] ;
   output [15:0]\FB_filter[1][0] ;
   output [15:0]\FB_filter[1][1] ;
   output [15:0]\FB_filter[1][2] ;
   output [15:0]\FB_filter[1][3] ;
   output [15:0]\FB_filter[1][4] ;
   output [15:0]\FB_filter[2][0] ;
   output [15:0]\FB_filter[2][1] ;
   output [15:0]\FB_filter[2][2] ;
   output [15:0]\FB_filter[2][3] ;
   output [15:0]\FB_filter[2][4] ;
   output [15:0]\FB_filter[3][0] ;
   output [15:0]\FB_filter[3][1] ;
   output [15:0]\FB_filter[3][2] ;
   output [15:0]\FB_filter[3][3] ;
   output [15:0]\FB_filter[3][4] ;
   output [15:0]\FB_filter[4][0] ;
   output [15:0]\FB_filter[4][1] ;
   output [15:0]\FB_filter[4][2] ;
   output [15:0]\FB_filter[4][3] ;
   output [15:0]\FB_filter[4][4] ;
   output [15:0]FB_index_filter;
   output [15:0]\FB_bias[0] ;
   output [15:0]\FB_bias[1] ;
   output [15:0]\FB_bias[2] ;
   output [15:0]\FB_bias[3] ;
   output [15:0]\FB_bias[4] ;
   output [15:0]\FB_bias[5] ;
   output [15:0]\FB_bias[6] ;
   output [15:0]\FB_bias[7] ;
   output [15:0]\FB_bias[8] ;
   output [15:0]\FB_bias[9] ;
   output [15:0]\FB_bias[10] ;
   output [15:0]\FB_bias[11] ;
   output [15:0]\FB_bias[12] ;
   output [15:0]\FB_bias[13] ;
   output [15:0]\FB_bias[14] ;
   output [15:0]\FB_bias[15] ;
   output [15:0]\FB_bias[16] ;
   output [15:0]\FB_bias[17] ;
   output [15:0]\FB_bias[18] ;
   output [15:0]\FB_bias[19] ;
   output [15:0]\FB_bias[20] ;
   output [15:0]\FB_bias[21] ;
   output [15:0]\FB_bias[22] ;
   output [15:0]\FB_bias[23] ;
   output [15:0]\FB_bias[24] ;
   output [15:0]\FB_bias[25] ;
   output [15:0]\FB_bias[26] ;
   output [15:0]\FB_bias[27] ;
   output [15:0]\FB_bias[28] ;
   output [15:0]\FB_bias[29] ;
   output [15:0]\FB_bias[30] ;
   output [15:0]\FB_bias[31] ;
   output [15:0]\FB_bias[32] ;
   output [15:0]\FB_bias[33] ;
   output [15:0]\FB_bias[34] ;
   output [15:0]\FB_bias[35] ;
   output [15:0]\FB_bias[36] ;
   output [15:0]\FB_bias[37] ;
   output [15:0]\FB_bias[38] ;
   output [15:0]\FB_bias[39] ;
   output [15:0]\FB_bias[40] ;
   output [15:0]\FB_bias[41] ;
   output [15:0]\FB_bias[42] ;
   output [15:0]\FB_bias[43] ;
   output [15:0]\FB_bias[44] ;
   output [15:0]\FB_bias[45] ;
   output [15:0]\FB_bias[46] ;
   output [15:0]\FB_bias[47] ;
   output [15:0]\FB_bias[48] ;
   output [15:0]\FB_bias[49] ;
   output [15:0]\FB_bias[50] ;
   output [15:0]\FB_bias[51] ;
   output [15:0]\FB_bias[52] ;
   output [15:0]\FB_bias[53] ;
   output [15:0]\FB_bias[54] ;
   output [15:0]\FB_bias[55] ;
   output [15:0]\FB_bias[56] ;
   output [15:0]\FB_bias[57] ;
   output [15:0]\FB_bias[58] ;
   output [15:0]\FB_bias[59] ;
   output [15:0]\FB_bias[60] ;
   output [15:0]\FB_bias[61] ;
   output [15:0]\FB_bias[62] ;
   output [15:0]\FB_bias[63] ;
   output [15:0]\FB_bias[64] ;
   output [15:0]\FB_bias[65] ;
   output [15:0]\FB_bias[66] ;
   output [15:0]\FB_bias[67] ;
   output [15:0]\FB_bias[68] ;
   output [15:0]\FB_bias[69] ;
   output [15:0]\FB_bias[70] ;
   output [15:0]\FB_bias[71] ;
   output [15:0]\FB_bias[72] ;
   output [15:0]\FB_bias[73] ;
   output [15:0]\FB_bias[74] ;
   output [15:0]\FB_bias[75] ;
   output [15:0]\FB_bias[76] ;
   output [15:0]\FB_bias[77] ;
   output [15:0]\FB_bias[78] ;
   output [15:0]\FB_bias[79] ;
   output [15:0]\FB_bias[80] ;
   output [15:0]\FB_bias[81] ;
   output [15:0]\FB_bias[82] ;
   output [15:0]\FB_bias[83] ;
   output [15:0]\FB_bias[84] ;
   output [15:0]\FB_bias[85] ;
   output [15:0]\FB_bias[86] ;
   output [15:0]\FB_bias[87] ;
   output [15:0]\FB_bias[88] ;
   output [15:0]\FB_bias[89] ;
   output [15:0]\FB_bias[90] ;
   output [15:0]\FB_bias[91] ;
   output [15:0]\FB_bias[92] ;
   output [15:0]\FB_bias[93] ;
   output [15:0]\FB_bias[94] ;
   output [15:0]\FB_bias[95] ;
   output [15:0]\FB_bias[96] ;
   output [15:0]\FB_bias[97] ;
   output [15:0]\FB_bias[98] ;
   output [15:0]\FB_bias[99] ;
   output [15:0]\FB_bias[100] ;
   output [15:0]\FB_bias[101] ;
   output [15:0]\FB_bias[102] ;
   output [15:0]\FB_bias[103] ;
   output [15:0]\FB_bias[104] ;
   output [15:0]\FB_bias[105] ;
   output [15:0]\FB_bias[106] ;
   output [15:0]\FB_bias[107] ;
   output [15:0]\FB_bias[108] ;
   output [15:0]\FB_bias[109] ;
   output [15:0]\FB_bias[110] ;
   output [15:0]\FB_bias[111] ;
   output [15:0]\FB_bias[112] ;
   output [15:0]\FB_bias[113] ;
   output [15:0]\FB_bias[114] ;
   output [15:0]\FB_bias[115] ;
   output [15:0]\FB_bias[116] ;
   output [15:0]\FB_bias[117] ;
   output [15:0]\FB_bias[118] ;
   output [15:0]\FB_bias[119] ;
   output FB_bias_or_filter;
   input FB_finish;

   wire n_2_2;
   wire n_2_4;
   wire n_2_5;
   wire n_2_6;
   wire n_2_7;
   wire n_2_8;
   wire n_2_9;
   wire n_2_10;
   wire n_2_11;
   wire n_2_12;
   wire n_2_13;
   wire n_2_14;
   wire n_2_15;
   wire n_2_16;
   wire n_2_17;
   wire n_2_0;
   wire n_2_1;
   wire n_2_3;
   wire n_2_0_0;
   wire n_2_0_1;
   wire n_2_0_2;
   wire n_2_0_3;
   wire n_0_0;
   wire n_0_1_0;
   wire n_0_1_1;
   wire n_0_16;
   wire n_0_15;
   wire n_0_14;
   wire n_0_13;
   wire n_0_12;
   wire n_0_11;
   wire n_0_10;
   wire n_0_9;
   wire n_0_8;
   wire n_0_7;
   wire n_0_6;
   wire n_0_5;
   wire n_0_4;
   wire n_0_3;
   wire n_0_2;
   wire n_0_1;

   DFF_X1 \RAM_address_reg[15]  (.D(n_2_1), .CK(n_2_2), .Q(n_0), .QN());
   DFF_X1 \RAM_address_reg[14]  (.D(n_2_0), .CK(n_2_2), .Q(n_1), .QN());
   DFF_X1 \RAM_address_reg[13]  (.D(n_2_17), .CK(n_2_2), .Q(n_2), .QN());
   DFF_X1 \RAM_address_reg[12]  (.D(n_2_16), .CK(n_2_2), .Q(n_3), .QN());
   DFF_X1 \RAM_address_reg[11]  (.D(n_2_15), .CK(n_2_2), .Q(n_4), .QN());
   DFF_X1 \RAM_address_reg[10]  (.D(n_2_14), .CK(n_2_2), .Q(n_5), .QN());
   DFF_X1 \RAM_address_reg[9]  (.D(n_2_13), .CK(n_2_2), .Q(n_6), .QN());
   DFF_X1 \RAM_address_reg[8]  (.D(n_2_12), .CK(n_2_2), .Q(n_7), .QN());
   DFF_X1 \RAM_address_reg[7]  (.D(n_2_11), .CK(n_2_2), .Q(n_8), .QN());
   DFF_X1 \RAM_address_reg[6]  (.D(n_2_10), .CK(n_2_2), .Q(n_9), .QN());
   DFF_X1 \RAM_address_reg[5]  (.D(n_2_9), .CK(n_2_2), .Q(n_10), .QN());
   DFF_X1 \RAM_address_reg[4]  (.D(n_2_8), .CK(n_2_2), .Q(n_11), .QN());
   DFF_X1 \RAM_address_reg[3]  (.D(n_2_7), .CK(n_2_2), .Q(n_12), .QN());
   DFF_X1 \RAM_address_reg[2]  (.D(n_2_6), .CK(n_2_2), .Q(n_13), .QN());
   DFF_X1 \RAM_address_reg[1]  (.D(n_2_5), .CK(n_2_2), .Q(n_14), .QN());
   DFF_X1 \RAM_address_reg[0]  (.D(n_2_4), .CK(n_2_2), .Q(n_15), .QN());
   CLKGATETST_X1 clk_gate_RAM_address_reg (.CK(clk), .E(n_2_3), .SE(1'b0), 
      .GCK(n_2_2));
   AND2_X1 i_2_0_0 (.A1(n_2_0_1), .A2(address[0]), .ZN(n_2_4));
   AND2_X1 i_2_0_1 (.A1(n_2_0_1), .A2(address[1]), .ZN(n_2_5));
   AND2_X1 i_2_0_2 (.A1(n_2_0_1), .A2(address[2]), .ZN(n_2_6));
   AND2_X1 i_2_0_3 (.A1(n_2_0_1), .A2(address[3]), .ZN(n_2_7));
   AND2_X1 i_2_0_4 (.A1(n_2_0_1), .A2(address[4]), .ZN(n_2_8));
   AND2_X1 i_2_0_5 (.A1(n_2_0_1), .A2(address[5]), .ZN(n_2_9));
   AND2_X1 i_2_0_6 (.A1(n_2_0_1), .A2(address[6]), .ZN(n_2_10));
   AND2_X1 i_2_0_7 (.A1(n_2_0_1), .A2(address[7]), .ZN(n_2_11));
   AND2_X1 i_2_0_8 (.A1(n_2_0_1), .A2(address[8]), .ZN(n_2_12));
   AND2_X1 i_2_0_9 (.A1(n_2_0_1), .A2(address[9]), .ZN(n_2_13));
   AND2_X1 i_2_0_10 (.A1(n_2_0_1), .A2(address[10]), .ZN(n_2_14));
   AND2_X1 i_2_0_11 (.A1(n_2_0_1), .A2(address[11]), .ZN(n_2_15));
   AND2_X1 i_2_0_12 (.A1(n_2_0_1), .A2(address[12]), .ZN(n_2_16));
   AND2_X1 i_2_0_13 (.A1(n_2_0_1), .A2(address[13]), .ZN(n_2_17));
   AND2_X1 i_2_0_14 (.A1(n_2_0_1), .A2(address[14]), .ZN(n_2_0));
   AND2_X1 i_2_0_15 (.A1(n_2_0_1), .A2(address[15]), .ZN(n_2_1));
   INV_X1 i_2_0_16 (.A(n_2_0_0), .ZN(n_2_3));
   OAI211_X1 i_2_0_17 (.A(start), .B(n_2_0_1), .C1(n_2_0_2), .C2(
      read_write_filter_bias[0]), .ZN(n_2_0_0));
   NAND2_X1 i_2_0_18 (.A1(n_2_0_3), .A2(read_write_filter_bias[0]), .ZN(n_2_0_1));
   OR4_X1 i_2_0_19 (.A1(filter_number[6]), .A2(n_2_0_3), .A3(filter_number[2]), 
      .A4(filter_number[10]), .ZN(n_2_0_2));
   INV_X1 i_2_0_20 (.A(read_write_filter_bias[1]), .ZN(n_2_0_3));
   DFF_X1 \RAM_address_reg[15]__0  (.D(n_0_16), .CK(n_0_0), .Q(n_0), .QN());
   DFF_X1 \RAM_address_reg[14]__0  (.D(n_0_15), .CK(n_0_0), .Q(n_1), .QN());
   DFF_X1 \RAM_address_reg[13]__0  (.D(n_0_14), .CK(n_0_0), .Q(n_2), .QN());
   DFF_X1 \RAM_address_reg[12]__0  (.D(n_0_13), .CK(n_0_0), .Q(n_3), .QN());
   DFF_X1 \RAM_address_reg[11]__0  (.D(n_0_12), .CK(n_0_0), .Q(n_4), .QN());
   DFF_X1 \RAM_address_reg[10]__0  (.D(n_0_11), .CK(n_0_0), .Q(n_5), .QN());
   DFF_X1 \RAM_address_reg[9]__0  (.D(n_0_10), .CK(n_0_0), .Q(n_6), .QN());
   DFF_X1 \RAM_address_reg[8]__0  (.D(n_0_9), .CK(n_0_0), .Q(n_7), .QN());
   DFF_X1 \RAM_address_reg[7]__0  (.D(n_0_8), .CK(n_0_0), .Q(n_8), .QN());
   DFF_X1 \RAM_address_reg[6]__0  (.D(n_0_7), .CK(n_0_0), .Q(n_9), .QN());
   DFF_X1 \RAM_address_reg[5]__0  (.D(n_0_6), .CK(n_0_0), .Q(n_10), .QN());
   DFF_X1 \RAM_address_reg[4]__0  (.D(n_0_5), .CK(n_0_0), .Q(n_11), .QN());
   DFF_X1 \RAM_address_reg[3]__0  (.D(n_0_4), .CK(n_0_0), .Q(n_12), .QN());
   DFF_X1 \RAM_address_reg[2]__0  (.D(n_0_3), .CK(n_0_0), .Q(n_13), .QN());
   DFF_X1 \RAM_address_reg[1]__0  (.D(n_0_2), .CK(n_0_0), .Q(n_14), .QN());
   DFF_X1 \RAM_address_reg[0]__0  (.D(n_0_1), .CK(n_0_0), .Q(n_15), .QN());
   INV_X1 i_0_0_0 (.A(clk), .ZN(n_0_0));
   NAND2_X1 i_0_1_0 (.A1(read_write_filter_bias[0]), .A2(start), .ZN(n_0_1_0));
   NOR2_X1 i_0_1_1 (.A1(n_0_1_0), .A2(read_write_filter_bias[1]), .ZN(n_0_1_1));
   MUX2_X1 i_0_1_2 (.A(n_0), .B(address[15]), .S(n_0_1_1), .Z(n_0_16));
   MUX2_X1 i_0_1_3 (.A(n_1), .B(address[14]), .S(n_0_1_1), .Z(n_0_15));
   MUX2_X1 i_0_1_4 (.A(n_2), .B(address[13]), .S(n_0_1_1), .Z(n_0_14));
   MUX2_X1 i_0_1_5 (.A(n_3), .B(address[12]), .S(n_0_1_1), .Z(n_0_13));
   MUX2_X1 i_0_1_6 (.A(n_4), .B(address[11]), .S(n_0_1_1), .Z(n_0_12));
   MUX2_X1 i_0_1_7 (.A(n_5), .B(address[10]), .S(n_0_1_1), .Z(n_0_11));
   MUX2_X1 i_0_1_8 (.A(n_6), .B(address[9]), .S(n_0_1_1), .Z(n_0_10));
   MUX2_X1 i_0_1_9 (.A(n_7), .B(address[8]), .S(n_0_1_1), .Z(n_0_9));
   MUX2_X1 i_0_1_10 (.A(n_8), .B(address[7]), .S(n_0_1_1), .Z(n_0_8));
   MUX2_X1 i_0_1_11 (.A(n_9), .B(address[6]), .S(n_0_1_1), .Z(n_0_7));
   MUX2_X1 i_0_1_12 (.A(n_10), .B(address[5]), .S(n_0_1_1), .Z(n_0_6));
   MUX2_X1 i_0_1_13 (.A(n_11), .B(address[4]), .S(n_0_1_1), .Z(n_0_5));
   MUX2_X1 i_0_1_14 (.A(n_12), .B(address[3]), .S(n_0_1_1), .Z(n_0_4));
   MUX2_X1 i_0_1_15 (.A(n_13), .B(address[2]), .S(n_0_1_1), .Z(n_0_3));
   MUX2_X1 i_0_1_16 (.A(n_14), .B(address[1]), .S(n_0_1_1), .Z(n_0_2));
   MUX2_X1 i_0_1_17 (.A(n_15), .B(address[0]), .S(n_0_1_1), .Z(n_0_1));
endmodule

module datapath__0_4270(p_0, p_1);
   input [15:0]p_0;
   output [15:0]p_1;

   HA_X1 i_1 (.A(p_0[1]), .B(p_0[0]), .CO(n_0), .S(p_1[1]));
   HA_X1 i_2 (.A(p_0[2]), .B(n_0), .CO(n_1), .S(p_1[2]));
   HA_X1 i_3 (.A(p_0[3]), .B(n_1), .CO(n_2), .S(p_1[3]));
   HA_X1 i_4 (.A(p_0[4]), .B(n_2), .CO(n_3), .S(p_1[4]));
   HA_X1 i_5 (.A(p_0[5]), .B(n_3), .CO(n_4), .S(p_1[5]));
   HA_X1 i_6 (.A(p_0[6]), .B(n_4), .CO(n_5), .S(p_1[6]));
   HA_X1 i_7 (.A(p_0[7]), .B(n_5), .CO(n_6), .S(p_1[7]));
   HA_X1 i_8 (.A(p_0[8]), .B(n_6), .CO(n_7), .S(p_1[8]));
   HA_X1 i_9 (.A(p_0[9]), .B(n_7), .CO(n_8), .S(p_1[9]));
   HA_X1 i_10 (.A(p_0[10]), .B(n_8), .CO(n_9), .S(p_1[10]));
   HA_X1 i_11 (.A(p_0[11]), .B(n_9), .CO(n_10), .S(p_1[11]));
   HA_X1 i_12 (.A(p_0[12]), .B(n_10), .CO(n_11), .S(p_1[12]));
   HA_X1 i_13 (.A(p_0[13]), .B(n_11), .CO(n_12), .S(p_1[13]));
   HA_X1 i_14 (.A(p_0[14]), .B(n_12), .CO(n_13), .S(p_1[14]));
   XOR2_X1 i_0 (.A(p_0[15]), .B(n_13), .Z(p_1[15]));
endmodule

module datapath__0_4273(p_0, p_1);
   input [15:0]p_0;
   output [15:0]p_1;

   HA_X1 i_1 (.A(p_0[1]), .B(p_0[0]), .CO(n_0), .S(p_1[1]));
   HA_X1 i_2 (.A(p_0[2]), .B(n_0), .CO(n_1), .S(p_1[2]));
   HA_X1 i_3 (.A(p_0[3]), .B(n_1), .CO(n_2), .S(p_1[3]));
   HA_X1 i_4 (.A(p_0[4]), .B(n_2), .CO(n_3), .S(p_1[4]));
   HA_X1 i_5 (.A(p_0[5]), .B(n_3), .CO(n_4), .S(p_1[5]));
   HA_X1 i_6 (.A(p_0[6]), .B(n_4), .CO(n_5), .S(p_1[6]));
   HA_X1 i_7 (.A(p_0[7]), .B(n_5), .CO(n_6), .S(p_1[7]));
   HA_X1 i_8 (.A(p_0[8]), .B(n_6), .CO(n_7), .S(p_1[8]));
   HA_X1 i_9 (.A(p_0[9]), .B(n_7), .CO(n_8), .S(p_1[9]));
   HA_X1 i_10 (.A(p_0[10]), .B(n_8), .CO(n_9), .S(p_1[10]));
   HA_X1 i_11 (.A(p_0[11]), .B(n_9), .CO(n_10), .S(p_1[11]));
   HA_X1 i_12 (.A(p_0[12]), .B(n_10), .CO(n_11), .S(p_1[12]));
   HA_X1 i_13 (.A(p_0[13]), .B(n_11), .CO(n_12), .S(p_1[13]));
   HA_X1 i_14 (.A(p_0[14]), .B(n_12), .CO(n_13), .S(p_1[14]));
   XOR2_X1 i_0 (.A(p_0[15]), .B(n_13), .Z(p_1[15]));
   INV_X1 i_15 (.A(p_0[0]), .ZN(p_1[0]));
endmodule

module datapath__0_4284(p_0, p_1);
   input [15:0]p_0;
   output [15:0]p_1;

   HA_X1 i_1 (.A(p_0[1]), .B(p_0[0]), .CO(n_0), .S(p_1[1]));
   HA_X1 i_2 (.A(p_0[2]), .B(n_0), .CO(n_1), .S(p_1[2]));
   HA_X1 i_3 (.A(p_0[3]), .B(n_1), .CO(n_2), .S(p_1[3]));
   HA_X1 i_4 (.A(p_0[4]), .B(n_2), .CO(n_3), .S(p_1[4]));
   HA_X1 i_5 (.A(p_0[5]), .B(n_3), .CO(n_4), .S(p_1[5]));
   HA_X1 i_6 (.A(p_0[6]), .B(n_4), .CO(n_5), .S(p_1[6]));
   HA_X1 i_7 (.A(p_0[7]), .B(n_5), .CO(n_6), .S(p_1[7]));
   HA_X1 i_8 (.A(p_0[8]), .B(n_6), .CO(n_7), .S(p_1[8]));
   HA_X1 i_9 (.A(p_0[9]), .B(n_7), .CO(n_8), .S(p_1[9]));
   HA_X1 i_10 (.A(p_0[10]), .B(n_8), .CO(n_9), .S(p_1[10]));
   HA_X1 i_11 (.A(p_0[11]), .B(n_9), .CO(n_10), .S(p_1[11]));
   HA_X1 i_12 (.A(p_0[12]), .B(n_10), .CO(n_11), .S(p_1[12]));
   HA_X1 i_13 (.A(p_0[13]), .B(n_11), .CO(n_12), .S(p_1[13]));
   HA_X1 i_14 (.A(p_0[14]), .B(n_12), .CO(n_13), .S(p_1[14]));
   XOR2_X1 i_0 (.A(p_0[15]), .B(n_13), .Z(p_1[15]));
   INV_X1 i_15 (.A(p_0[0]), .ZN(p_1[0]));
endmodule

module datapath__0_4288(featureMapSize, p_0, p_1);
   input [6:0]featureMapSize;
   input [15:0]p_0;
   output [15:0]p_1;

   HA_X1 i_0 (.A(featureMapSize[0]), .B(p_0[0]), .CO(n_0), .S(p_1[0]));
   FA_X1 i_1 (.A(featureMapSize[1]), .B(p_0[1]), .CI(n_0), .CO(n_1), .S(p_1[1]));
   FA_X1 i_2 (.A(featureMapSize[2]), .B(p_0[2]), .CI(n_1), .CO(n_2), .S(p_1[2]));
   FA_X1 i_3 (.A(featureMapSize[3]), .B(p_0[3]), .CI(n_2), .CO(n_3), .S(p_1[3]));
   FA_X1 i_4 (.A(featureMapSize[4]), .B(p_0[4]), .CI(n_3), .CO(n_4), .S(p_1[4]));
   FA_X1 i_5 (.A(featureMapSize[5]), .B(p_0[5]), .CI(n_4), .CO(n_5), .S(p_1[5]));
   HA_X1 i_6 (.A(p_0[6]), .B(n_5), .CO(n_6), .S(p_1[6]));
   HA_X1 i_7 (.A(p_0[7]), .B(n_6), .CO(n_7), .S(p_1[7]));
   HA_X1 i_8 (.A(p_0[8]), .B(n_7), .CO(n_8), .S(p_1[8]));
   HA_X1 i_9 (.A(p_0[9]), .B(n_8), .CO(n_9), .S(p_1[9]));
   HA_X1 i_10 (.A(p_0[10]), .B(n_9), .CO(n_10), .S(p_1[10]));
   HA_X1 i_11 (.A(p_0[11]), .B(n_10), .CO(n_11), .S(p_1[11]));
   HA_X1 i_12 (.A(p_0[12]), .B(n_11), .CO(n_12), .S(p_1[12]));
   HA_X1 i_13 (.A(p_0[13]), .B(n_12), .CO(n_13), .S(p_1[13]));
   HA_X1 i_14 (.A(p_0[14]), .B(n_13), .CO(n_14), .S(p_1[14]));
   XOR2_X1 i_15 (.A(p_0[15]), .B(n_14), .Z(p_1[15]));
endmodule

module datapath__0_4294(p_0, p_1, p_2);
   input [10:0]p_0;
   input [15:0]p_1;
   output [15:0]p_2;

   FA_X1 i_26 (.A(p_1[2]), .B(n_0), .CI(n_23), .CO(n_24), .S(p_2[2]));
   FA_X1 i_27 (.A(n_1), .B(n_2), .CI(n_24), .CO(n_25), .S(p_2[3]));
   FA_X1 i_28 (.A(n_3), .B(n_4), .CI(n_25), .CO(n_26), .S(p_2[4]));
   FA_X1 i_29 (.A(n_5), .B(n_6), .CI(n_26), .CO(n_27), .S(p_2[5]));
   FA_X1 i_30 (.A(n_7), .B(n_8), .CI(n_27), .CO(n_28), .S(p_2[6]));
   FA_X1 i_31 (.A(n_9), .B(n_10), .CI(n_28), .CO(n_29), .S(p_2[7]));
   FA_X1 i_32 (.A(n_11), .B(n_12), .CI(n_29), .CO(n_30), .S(p_2[8]));
   FA_X1 i_33 (.A(n_13), .B(n_14), .CI(n_30), .CO(n_31), .S(p_2[9]));
   FA_X1 i_34 (.A(n_15), .B(n_16), .CI(n_31), .CO(n_32), .S(p_2[10]));
   FA_X1 i_35 (.A(n_17), .B(n_19), .CI(n_32), .CO(n_33), .S(p_2[11]));
   FA_X1 i_36 (.A(p_1[12]), .B(n_19), .CI(n_33), .CO(n_34), .S(p_2[12]));
   FA_X1 i_37 (.A(p_1[13]), .B(n_19), .CI(n_34), .CO(n_35), .S(p_2[13]));
   FA_X1 i_38 (.A(p_1[14]), .B(n_19), .CI(n_35), .CO(n_36), .S(p_2[14]));
   XNOR2_X1 i_0 (.A(p_0[10]), .B(p_1[10]), .ZN(n_16));
   NOR2_X1 i_1 (.A1(n_22), .A2(p_0[10]), .ZN(n_17));
   OR2_X1 i_2 (.A1(p_0[9]), .A2(p_1[9]), .ZN(n_15));
   XNOR2_X1 i_3 (.A(p_0[9]), .B(p_1[9]), .ZN(n_14));
   OR2_X1 i_4 (.A1(p_0[8]), .A2(p_1[8]), .ZN(n_13));
   XNOR2_X1 i_5 (.A(p_0[8]), .B(p_1[8]), .ZN(n_12));
   OR2_X1 i_6 (.A1(p_0[7]), .A2(p_1[7]), .ZN(n_11));
   XNOR2_X1 i_7 (.A(p_0[7]), .B(p_1[7]), .ZN(n_10));
   OR2_X1 i_8 (.A1(p_0[6]), .A2(p_1[6]), .ZN(n_9));
   XNOR2_X1 i_9 (.A(p_0[6]), .B(p_1[6]), .ZN(n_8));
   OR2_X1 i_10 (.A1(p_0[5]), .A2(p_1[5]), .ZN(n_7));
   XNOR2_X1 i_11 (.A(p_0[5]), .B(p_1[5]), .ZN(n_6));
   OR2_X1 i_12 (.A1(p_0[4]), .A2(p_1[4]), .ZN(n_5));
   XNOR2_X1 i_13 (.A(p_0[4]), .B(p_1[4]), .ZN(n_4));
   OR2_X1 i_14 (.A1(p_0[3]), .A2(p_1[3]), .ZN(n_3));
   XNOR2_X1 i_15 (.A(p_0[3]), .B(p_1[3]), .ZN(n_2));
   OR2_X1 i_16 (.A1(p_0[2]), .A2(p_0[0]), .ZN(n_1));
   XNOR2_X1 i_17 (.A(p_0[2]), .B(p_0[0]), .ZN(n_0));
   XNOR2_X1 i_18 (.A(p_0[0]), .B(n_21), .ZN(p_2[0]));
   XNOR2_X1 i_19 (.A(p_1[1]), .B(n_18), .ZN(p_2[1]));
   OR2_X1 i_20 (.A1(n_18), .A2(p_1[1]), .ZN(n_23));
   NAND2_X1 i_21 (.A1(n_21), .A2(p_0[0]), .ZN(n_18));
   XNOR2_X1 i_22 (.A(p_1[15]), .B(n_20), .ZN(p_2[15]));
   XNOR2_X1 i_23 (.A(n_19), .B(n_36), .ZN(n_20));
   INV_X1 i_24 (.A(p_1[0]), .ZN(n_21));
   INV_X1 i_25 (.A(p_1[10]), .ZN(n_22));
   INV_X1 i_39 (.A(p_1[11]), .ZN(n_19));
endmodule

module datapath__0_4295(p_0, p_1, p_2);
   input [11:0]p_0;
   input [15:0]p_1;
   output [15:0]p_2;

   INV_X1 i_1 (.A(p_1[12]), .ZN(n_1));
   HA_X1 i_2 (.A(p_0[0]), .B(p_1[0]), .CO(n_2), .S(p_2[0]));
   HA_X1 i_3 (.A(p_1[1]), .B(n_2), .CO(n_3), .S(p_2[1]));
   FA_X1 i_4 (.A(p_0[2]), .B(p_1[2]), .CI(n_3), .CO(n_4), .S(p_2[2]));
   FA_X1 i_5 (.A(p_0[3]), .B(p_1[3]), .CI(n_4), .CO(n_5), .S(p_2[3]));
   FA_X1 i_6 (.A(p_0[4]), .B(p_1[4]), .CI(n_5), .CO(n_6), .S(p_2[4]));
   FA_X1 i_7 (.A(p_0[5]), .B(p_1[5]), .CI(n_6), .CO(n_7), .S(p_2[5]));
   FA_X1 i_8 (.A(p_0[6]), .B(p_1[6]), .CI(n_7), .CO(n_8), .S(p_2[6]));
   FA_X1 i_9 (.A(p_0[7]), .B(p_1[7]), .CI(n_8), .CO(n_9), .S(p_2[7]));
   FA_X1 i_10 (.A(p_0[8]), .B(p_1[8]), .CI(n_9), .CO(n_10), .S(p_2[8]));
   FA_X1 i_11 (.A(p_0[9]), .B(p_1[9]), .CI(n_10), .CO(n_11), .S(p_2[9]));
   FA_X1 i_12 (.A(p_0[10]), .B(p_1[10]), .CI(n_11), .CO(n_12), .S(p_2[10]));
   FA_X1 i_13 (.A(p_1[11]), .B(1'b0), .CI(n_12), .CO(n_13), .S(p_2[11]));
   FA_X1 i_14 (.A(1'b1), .B(n_1), .CI(n_13), .CO(n_14), .S(p_2[12]));
   FA_X1 i_15 (.A(p_1[13]), .B(n_1), .CI(n_14), .CO(n_15), .S(p_2[13]));
   FA_X1 i_16 (.A(p_1[14]), .B(n_1), .CI(n_15), .CO(n_16), .S(p_2[14]));
   XNOR2_X1 i_17 (.A(p_1[15]), .B(n_1), .ZN(n_0));
   XNOR2_X1 i_18 (.A(n_0), .B(n_16), .ZN(p_2[15]));
endmodule

module datapath__0_4312(filterCounter, p_0);
   input [31:0]filterCounter;
   output [31:0]p_0;

   HA_X1 i_1 (.A(filterCounter[1]), .B(filterCounter[0]), .CO(n_0), .S(p_0[1]));
   HA_X1 i_2 (.A(filterCounter[2]), .B(n_0), .CO(n_1), .S(p_0[2]));
   HA_X1 i_3 (.A(filterCounter[3]), .B(n_1), .CO(n_2), .S(p_0[3]));
   HA_X1 i_4 (.A(filterCounter[4]), .B(n_2), .CO(n_3), .S(p_0[4]));
   HA_X1 i_5 (.A(filterCounter[5]), .B(n_3), .CO(n_4), .S(p_0[5]));
   HA_X1 i_6 (.A(filterCounter[6]), .B(n_4), .CO(n_5), .S(p_0[6]));
   HA_X1 i_7 (.A(filterCounter[7]), .B(n_5), .CO(n_6), .S(p_0[7]));
   HA_X1 i_8 (.A(filterCounter[8]), .B(n_6), .CO(n_7), .S(p_0[8]));
   HA_X1 i_9 (.A(filterCounter[9]), .B(n_7), .CO(n_8), .S(p_0[9]));
   HA_X1 i_10 (.A(filterCounter[10]), .B(n_8), .CO(n_9), .S(p_0[10]));
   HA_X1 i_11 (.A(filterCounter[11]), .B(n_9), .CO(n_10), .S(p_0[11]));
   HA_X1 i_12 (.A(filterCounter[12]), .B(n_10), .CO(n_11), .S(p_0[12]));
   HA_X1 i_13 (.A(filterCounter[13]), .B(n_11), .CO(n_12), .S(p_0[13]));
   HA_X1 i_14 (.A(filterCounter[14]), .B(n_12), .CO(n_13), .S(p_0[14]));
   HA_X1 i_15 (.A(filterCounter[15]), .B(n_13), .CO(n_14), .S(p_0[15]));
   HA_X1 i_16 (.A(filterCounter[16]), .B(n_14), .CO(n_15), .S(p_0[16]));
   HA_X1 i_17 (.A(filterCounter[17]), .B(n_15), .CO(n_16), .S(p_0[17]));
   HA_X1 i_18 (.A(filterCounter[18]), .B(n_16), .CO(n_17), .S(p_0[18]));
   HA_X1 i_19 (.A(filterCounter[19]), .B(n_17), .CO(n_18), .S(p_0[19]));
   HA_X1 i_20 (.A(filterCounter[20]), .B(n_18), .CO(n_19), .S(p_0[20]));
   HA_X1 i_21 (.A(filterCounter[21]), .B(n_19), .CO(n_20), .S(p_0[21]));
   HA_X1 i_22 (.A(filterCounter[22]), .B(n_20), .CO(n_21), .S(p_0[22]));
   HA_X1 i_23 (.A(filterCounter[23]), .B(n_21), .CO(n_22), .S(p_0[23]));
   HA_X1 i_24 (.A(filterCounter[24]), .B(n_22), .CO(n_23), .S(p_0[24]));
   HA_X1 i_25 (.A(filterCounter[25]), .B(n_23), .CO(n_24), .S(p_0[25]));
   HA_X1 i_26 (.A(filterCounter[26]), .B(n_24), .CO(n_25), .S(p_0[26]));
   HA_X1 i_27 (.A(filterCounter[27]), .B(n_25), .CO(n_26), .S(p_0[27]));
   HA_X1 i_28 (.A(filterCounter[28]), .B(n_26), .CO(n_27), .S(p_0[28]));
   HA_X1 i_29 (.A(filterCounter[29]), .B(n_27), .CO(n_28), .S(p_0[29]));
   HA_X1 i_30 (.A(filterCounter[30]), .B(n_28), .CO(n_29), .S(p_0[30]));
   XOR2_X1 i_0 (.A(filterCounter[31]), .B(n_29), .Z(p_0[31]));
endmodule

module datapath__0_4318(convWindowX, p_0);
   input [31:0]convWindowX;
   output [31:0]p_0;

   HA_X1 i_1 (.A(convWindowX[1]), .B(convWindowX[0]), .CO(n_0), .S(p_0[1]));
   HA_X1 i_2 (.A(convWindowX[2]), .B(n_0), .CO(n_1), .S(p_0[2]));
   HA_X1 i_3 (.A(convWindowX[3]), .B(n_1), .CO(n_2), .S(p_0[3]));
   HA_X1 i_4 (.A(convWindowX[4]), .B(n_2), .CO(n_3), .S(p_0[4]));
   HA_X1 i_5 (.A(convWindowX[5]), .B(n_3), .CO(n_4), .S(p_0[5]));
   HA_X1 i_6 (.A(convWindowX[6]), .B(n_4), .CO(n_5), .S(p_0[6]));
   HA_X1 i_7 (.A(convWindowX[7]), .B(n_5), .CO(n_6), .S(p_0[7]));
   HA_X1 i_8 (.A(convWindowX[8]), .B(n_6), .CO(n_7), .S(p_0[8]));
   HA_X1 i_9 (.A(convWindowX[9]), .B(n_7), .CO(n_8), .S(p_0[9]));
   HA_X1 i_10 (.A(convWindowX[10]), .B(n_8), .CO(n_9), .S(p_0[10]));
   HA_X1 i_11 (.A(convWindowX[11]), .B(n_9), .CO(n_10), .S(p_0[11]));
   HA_X1 i_12 (.A(convWindowX[12]), .B(n_10), .CO(n_11), .S(p_0[12]));
   HA_X1 i_13 (.A(convWindowX[13]), .B(n_11), .CO(n_12), .S(p_0[13]));
   HA_X1 i_14 (.A(convWindowX[14]), .B(n_12), .CO(n_13), .S(p_0[14]));
   HA_X1 i_15 (.A(convWindowX[15]), .B(n_13), .CO(n_14), .S(p_0[15]));
   HA_X1 i_16 (.A(convWindowX[16]), .B(n_14), .CO(n_15), .S(p_0[16]));
   HA_X1 i_17 (.A(convWindowX[17]), .B(n_15), .CO(n_16), .S(p_0[17]));
   HA_X1 i_18 (.A(convWindowX[18]), .B(n_16), .CO(n_17), .S(p_0[18]));
   HA_X1 i_19 (.A(convWindowX[19]), .B(n_17), .CO(n_18), .S(p_0[19]));
   HA_X1 i_20 (.A(convWindowX[20]), .B(n_18), .CO(n_19), .S(p_0[20]));
   HA_X1 i_21 (.A(convWindowX[21]), .B(n_19), .CO(n_20), .S(p_0[21]));
   HA_X1 i_22 (.A(convWindowX[22]), .B(n_20), .CO(n_21), .S(p_0[22]));
   HA_X1 i_23 (.A(convWindowX[23]), .B(n_21), .CO(n_22), .S(p_0[23]));
   HA_X1 i_24 (.A(convWindowX[24]), .B(n_22), .CO(n_23), .S(p_0[24]));
   HA_X1 i_25 (.A(convWindowX[25]), .B(n_23), .CO(n_24), .S(p_0[25]));
   HA_X1 i_26 (.A(convWindowX[26]), .B(n_24), .CO(n_25), .S(p_0[26]));
   HA_X1 i_27 (.A(convWindowX[27]), .B(n_25), .CO(n_26), .S(p_0[27]));
   HA_X1 i_28 (.A(convWindowX[28]), .B(n_26), .CO(n_27), .S(p_0[28]));
   HA_X1 i_29 (.A(convWindowX[29]), .B(n_27), .CO(n_28), .S(p_0[29]));
   HA_X1 i_30 (.A(convWindowX[30]), .B(n_28), .CO(n_29), .S(p_0[30]));
   XOR2_X1 i_0 (.A(convWindowX[31]), .B(n_29), .Z(p_0[31]));
endmodule

module datapath__0_4321(kernelCounter, p_0);
   input [31:0]kernelCounter;
   output [31:0]p_0;

   HA_X1 i_1 (.A(kernelCounter[1]), .B(kernelCounter[0]), .CO(n_0), .S(p_0[1]));
   HA_X1 i_2 (.A(kernelCounter[2]), .B(n_0), .CO(n_1), .S(p_0[2]));
   HA_X1 i_3 (.A(kernelCounter[3]), .B(n_1), .CO(n_2), .S(p_0[3]));
   HA_X1 i_4 (.A(kernelCounter[4]), .B(n_2), .CO(n_3), .S(p_0[4]));
   HA_X1 i_5 (.A(kernelCounter[5]), .B(n_3), .CO(n_4), .S(p_0[5]));
   HA_X1 i_6 (.A(kernelCounter[6]), .B(n_4), .CO(n_5), .S(p_0[6]));
   HA_X1 i_7 (.A(kernelCounter[7]), .B(n_5), .CO(n_6), .S(p_0[7]));
   HA_X1 i_8 (.A(kernelCounter[8]), .B(n_6), .CO(n_7), .S(p_0[8]));
   HA_X1 i_9 (.A(kernelCounter[9]), .B(n_7), .CO(n_8), .S(p_0[9]));
   HA_X1 i_10 (.A(kernelCounter[10]), .B(n_8), .CO(n_9), .S(p_0[10]));
   HA_X1 i_11 (.A(kernelCounter[11]), .B(n_9), .CO(n_10), .S(p_0[11]));
   HA_X1 i_12 (.A(kernelCounter[12]), .B(n_10), .CO(n_11), .S(p_0[12]));
   HA_X1 i_13 (.A(kernelCounter[13]), .B(n_11), .CO(n_12), .S(p_0[13]));
   HA_X1 i_14 (.A(kernelCounter[14]), .B(n_12), .CO(n_13), .S(p_0[14]));
   HA_X1 i_15 (.A(kernelCounter[15]), .B(n_13), .CO(n_14), .S(p_0[15]));
   HA_X1 i_16 (.A(kernelCounter[16]), .B(n_14), .CO(n_15), .S(p_0[16]));
   HA_X1 i_17 (.A(kernelCounter[17]), .B(n_15), .CO(n_16), .S(p_0[17]));
   HA_X1 i_18 (.A(kernelCounter[18]), .B(n_16), .CO(n_17), .S(p_0[18]));
   HA_X1 i_19 (.A(kernelCounter[19]), .B(n_17), .CO(n_18), .S(p_0[19]));
   HA_X1 i_20 (.A(kernelCounter[20]), .B(n_18), .CO(n_19), .S(p_0[20]));
   HA_X1 i_21 (.A(kernelCounter[21]), .B(n_19), .CO(n_20), .S(p_0[21]));
   HA_X1 i_22 (.A(kernelCounter[22]), .B(n_20), .CO(n_21), .S(p_0[22]));
   HA_X1 i_23 (.A(kernelCounter[23]), .B(n_21), .CO(n_22), .S(p_0[23]));
   HA_X1 i_24 (.A(kernelCounter[24]), .B(n_22), .CO(n_23), .S(p_0[24]));
   HA_X1 i_25 (.A(kernelCounter[25]), .B(n_23), .CO(n_24), .S(p_0[25]));
   HA_X1 i_26 (.A(kernelCounter[26]), .B(n_24), .CO(n_25), .S(p_0[26]));
   HA_X1 i_27 (.A(kernelCounter[27]), .B(n_25), .CO(n_26), .S(p_0[27]));
   HA_X1 i_28 (.A(kernelCounter[28]), .B(n_26), .CO(n_27), .S(p_0[28]));
   HA_X1 i_29 (.A(kernelCounter[29]), .B(n_27), .CO(n_28), .S(p_0[29]));
   HA_X1 i_30 (.A(kernelCounter[30]), .B(n_28), .CO(n_29), .S(p_0[30]));
   XOR2_X1 i_0 (.A(kernelCounter[31]), .B(n_29), .Z(p_0[31]));
   INV_X1 i_31 (.A(kernelCounter[0]), .ZN(p_0[0]));
endmodule

module datapath__0_4332(poolingWindowY, p_0);
   input [31:0]poolingWindowY;
   output [31:0]p_0;

   HA_X1 i_1 (.A(poolingWindowY[2]), .B(poolingWindowY[1]), .CO(n_0), .S(p_0[2]));
   HA_X1 i_2 (.A(poolingWindowY[3]), .B(n_0), .CO(n_1), .S(p_0[3]));
   HA_X1 i_3 (.A(poolingWindowY[4]), .B(n_1), .CO(n_2), .S(p_0[4]));
   HA_X1 i_4 (.A(poolingWindowY[5]), .B(n_2), .CO(n_3), .S(p_0[5]));
   HA_X1 i_5 (.A(poolingWindowY[6]), .B(n_3), .CO(n_4), .S(p_0[6]));
   HA_X1 i_6 (.A(poolingWindowY[7]), .B(n_4), .CO(n_5), .S(p_0[7]));
   HA_X1 i_7 (.A(poolingWindowY[8]), .B(n_5), .CO(n_6), .S(p_0[8]));
   HA_X1 i_8 (.A(poolingWindowY[9]), .B(n_6), .CO(n_7), .S(p_0[9]));
   HA_X1 i_9 (.A(poolingWindowY[10]), .B(n_7), .CO(n_8), .S(p_0[10]));
   HA_X1 i_10 (.A(poolingWindowY[11]), .B(n_8), .CO(n_9), .S(p_0[11]));
   HA_X1 i_11 (.A(poolingWindowY[12]), .B(n_9), .CO(n_10), .S(p_0[12]));
   HA_X1 i_12 (.A(poolingWindowY[13]), .B(n_10), .CO(n_11), .S(p_0[13]));
   HA_X1 i_13 (.A(poolingWindowY[14]), .B(n_11), .CO(n_12), .S(p_0[14]));
   HA_X1 i_14 (.A(poolingWindowY[15]), .B(n_12), .CO(n_13), .S(p_0[15]));
   HA_X1 i_15 (.A(poolingWindowY[16]), .B(n_13), .CO(n_14), .S(p_0[16]));
   HA_X1 i_16 (.A(poolingWindowY[17]), .B(n_14), .CO(n_15), .S(p_0[17]));
   HA_X1 i_17 (.A(poolingWindowY[18]), .B(n_15), .CO(n_16), .S(p_0[18]));
   HA_X1 i_18 (.A(poolingWindowY[19]), .B(n_16), .CO(n_17), .S(p_0[19]));
   HA_X1 i_19 (.A(poolingWindowY[20]), .B(n_17), .CO(n_18), .S(p_0[20]));
   HA_X1 i_20 (.A(poolingWindowY[21]), .B(n_18), .CO(n_19), .S(p_0[21]));
   HA_X1 i_21 (.A(poolingWindowY[22]), .B(n_19), .CO(n_20), .S(p_0[22]));
   HA_X1 i_22 (.A(poolingWindowY[23]), .B(n_20), .CO(n_21), .S(p_0[23]));
   HA_X1 i_23 (.A(poolingWindowY[24]), .B(n_21), .CO(n_22), .S(p_0[24]));
   HA_X1 i_24 (.A(poolingWindowY[25]), .B(n_22), .CO(n_23), .S(p_0[25]));
   HA_X1 i_25 (.A(poolingWindowY[26]), .B(n_23), .CO(n_24), .S(p_0[26]));
   HA_X1 i_26 (.A(poolingWindowY[27]), .B(n_24), .CO(n_25), .S(p_0[27]));
   HA_X1 i_27 (.A(poolingWindowY[28]), .B(n_25), .CO(n_26), .S(p_0[28]));
   HA_X1 i_28 (.A(poolingWindowY[29]), .B(n_26), .CO(n_27), .S(p_0[29]));
   HA_X1 i_29 (.A(poolingWindowY[30]), .B(n_27), .CO(n_28), .S(p_0[30]));
   XOR2_X1 i_0 (.A(poolingWindowY[31]), .B(n_28), .Z(p_0[31]));
   INV_X1 i_30 (.A(poolingWindowY[1]), .ZN(p_0[1]));
endmodule

module datapath__0_4335(poolingWindowX, p_0);
   input [31:0]poolingWindowX;
   output [31:0]p_0;

   HA_X1 i_1 (.A(poolingWindowX[2]), .B(poolingWindowX[1]), .CO(n_0), .S(p_0[2]));
   HA_X1 i_2 (.A(poolingWindowX[3]), .B(n_0), .CO(n_1), .S(p_0[3]));
   HA_X1 i_3 (.A(poolingWindowX[4]), .B(n_1), .CO(n_2), .S(p_0[4]));
   HA_X1 i_4 (.A(poolingWindowX[5]), .B(n_2), .CO(n_3), .S(p_0[5]));
   HA_X1 i_5 (.A(poolingWindowX[6]), .B(n_3), .CO(n_4), .S(p_0[6]));
   HA_X1 i_6 (.A(poolingWindowX[7]), .B(n_4), .CO(n_5), .S(p_0[7]));
   HA_X1 i_7 (.A(poolingWindowX[8]), .B(n_5), .CO(n_6), .S(p_0[8]));
   HA_X1 i_8 (.A(poolingWindowX[9]), .B(n_6), .CO(n_7), .S(p_0[9]));
   HA_X1 i_9 (.A(poolingWindowX[10]), .B(n_7), .CO(n_8), .S(p_0[10]));
   HA_X1 i_10 (.A(poolingWindowX[11]), .B(n_8), .CO(n_9), .S(p_0[11]));
   HA_X1 i_11 (.A(poolingWindowX[12]), .B(n_9), .CO(n_10), .S(p_0[12]));
   HA_X1 i_12 (.A(poolingWindowX[13]), .B(n_10), .CO(n_11), .S(p_0[13]));
   HA_X1 i_13 (.A(poolingWindowX[14]), .B(n_11), .CO(n_12), .S(p_0[14]));
   HA_X1 i_14 (.A(poolingWindowX[15]), .B(n_12), .CO(n_13), .S(p_0[15]));
   HA_X1 i_15 (.A(poolingWindowX[16]), .B(n_13), .CO(n_14), .S(p_0[16]));
   HA_X1 i_16 (.A(poolingWindowX[17]), .B(n_14), .CO(n_15), .S(p_0[17]));
   HA_X1 i_17 (.A(poolingWindowX[18]), .B(n_15), .CO(n_16), .S(p_0[18]));
   HA_X1 i_18 (.A(poolingWindowX[19]), .B(n_16), .CO(n_17), .S(p_0[19]));
   HA_X1 i_19 (.A(poolingWindowX[20]), .B(n_17), .CO(n_18), .S(p_0[20]));
   HA_X1 i_20 (.A(poolingWindowX[21]), .B(n_18), .CO(n_19), .S(p_0[21]));
   HA_X1 i_21 (.A(poolingWindowX[22]), .B(n_19), .CO(n_20), .S(p_0[22]));
   HA_X1 i_22 (.A(poolingWindowX[23]), .B(n_20), .CO(n_21), .S(p_0[23]));
   HA_X1 i_23 (.A(poolingWindowX[24]), .B(n_21), .CO(n_22), .S(p_0[24]));
   HA_X1 i_24 (.A(poolingWindowX[25]), .B(n_22), .CO(n_23), .S(p_0[25]));
   HA_X1 i_25 (.A(poolingWindowX[26]), .B(n_23), .CO(n_24), .S(p_0[26]));
   HA_X1 i_26 (.A(poolingWindowX[27]), .B(n_24), .CO(n_25), .S(p_0[27]));
   HA_X1 i_27 (.A(poolingWindowX[28]), .B(n_25), .CO(n_26), .S(p_0[28]));
   HA_X1 i_28 (.A(poolingWindowX[29]), .B(n_26), .CO(n_27), .S(p_0[29]));
   HA_X1 i_29 (.A(poolingWindowX[30]), .B(n_27), .CO(n_28), .S(p_0[30]));
   XOR2_X1 i_0 (.A(poolingWindowX[31]), .B(n_28), .Z(p_0[31]));
   INV_X1 i_30 (.A(poolingWindowX[1]), .ZN(p_0[1]));
endmodule

module datapath__0_4338(poolingCounter, p_0);
   input [31:0]poolingCounter;
   output [31:0]p_0;

   HA_X1 i_1 (.A(poolingCounter[1]), .B(poolingCounter[0]), .CO(n_0), .S(p_0[1]));
   HA_X1 i_2 (.A(poolingCounter[2]), .B(n_0), .CO(n_1), .S(p_0[2]));
   HA_X1 i_3 (.A(poolingCounter[3]), .B(n_1), .CO(n_2), .S(p_0[3]));
   HA_X1 i_4 (.A(poolingCounter[4]), .B(n_2), .CO(n_3), .S(p_0[4]));
   HA_X1 i_5 (.A(poolingCounter[5]), .B(n_3), .CO(n_4), .S(p_0[5]));
   HA_X1 i_6 (.A(poolingCounter[6]), .B(n_4), .CO(n_5), .S(p_0[6]));
   HA_X1 i_7 (.A(poolingCounter[7]), .B(n_5), .CO(n_6), .S(p_0[7]));
   HA_X1 i_8 (.A(poolingCounter[8]), .B(n_6), .CO(n_7), .S(p_0[8]));
   HA_X1 i_9 (.A(poolingCounter[9]), .B(n_7), .CO(n_8), .S(p_0[9]));
   HA_X1 i_10 (.A(poolingCounter[10]), .B(n_8), .CO(n_9), .S(p_0[10]));
   HA_X1 i_11 (.A(poolingCounter[11]), .B(n_9), .CO(n_10), .S(p_0[11]));
   HA_X1 i_12 (.A(poolingCounter[12]), .B(n_10), .CO(n_11), .S(p_0[12]));
   HA_X1 i_13 (.A(poolingCounter[13]), .B(n_11), .CO(n_12), .S(p_0[13]));
   HA_X1 i_14 (.A(poolingCounter[14]), .B(n_12), .CO(n_13), .S(p_0[14]));
   HA_X1 i_15 (.A(poolingCounter[15]), .B(n_13), .CO(n_14), .S(p_0[15]));
   HA_X1 i_16 (.A(poolingCounter[16]), .B(n_14), .CO(n_15), .S(p_0[16]));
   HA_X1 i_17 (.A(poolingCounter[17]), .B(n_15), .CO(n_16), .S(p_0[17]));
   HA_X1 i_18 (.A(poolingCounter[18]), .B(n_16), .CO(n_17), .S(p_0[18]));
   HA_X1 i_19 (.A(poolingCounter[19]), .B(n_17), .CO(n_18), .S(p_0[19]));
   HA_X1 i_20 (.A(poolingCounter[20]), .B(n_18), .CO(n_19), .S(p_0[20]));
   HA_X1 i_21 (.A(poolingCounter[21]), .B(n_19), .CO(n_20), .S(p_0[21]));
   HA_X1 i_22 (.A(poolingCounter[22]), .B(n_20), .CO(n_21), .S(p_0[22]));
   HA_X1 i_23 (.A(poolingCounter[23]), .B(n_21), .CO(n_22), .S(p_0[23]));
   HA_X1 i_24 (.A(poolingCounter[24]), .B(n_22), .CO(n_23), .S(p_0[24]));
   HA_X1 i_25 (.A(poolingCounter[25]), .B(n_23), .CO(n_24), .S(p_0[25]));
   HA_X1 i_26 (.A(poolingCounter[26]), .B(n_24), .CO(n_25), .S(p_0[26]));
   HA_X1 i_27 (.A(poolingCounter[27]), .B(n_25), .CO(n_26), .S(p_0[27]));
   HA_X1 i_28 (.A(poolingCounter[28]), .B(n_26), .CO(n_27), .S(p_0[28]));
   HA_X1 i_29 (.A(poolingCounter[29]), .B(n_27), .CO(n_28), .S(p_0[29]));
   HA_X1 i_30 (.A(poolingCounter[30]), .B(n_28), .CO(n_29), .S(p_0[30]));
   XOR2_X1 i_0 (.A(poolingCounter[31]), .B(n_29), .Z(p_0[31]));
endmodule

module CNN(start, reset, finish, clk, \filter[0][0] , \filter[0][1] , 
      \filter[0][2] , \filter[0][3] , \filter[0][4] , \filter[1][0] , 
      \filter[1][1] , \filter[1][2] , \filter[1][3] , \filter[1][4] , 
      \filter[2][0] , \filter[2][1] , \filter[2][2] , \filter[2][3] , 
      \filter[2][4] , \filter[3][0] , \filter[3][1] , \filter[3][2] , 
      \filter[3][3] , \filter[3][4] , \filter[4][0] , \filter[4][1] , 
      \filter[4][2] , \filter[4][3] , \filter[4][4] , FB_index_bias, 
      FB_output_bias, index_filter, DMA_start, DMA_finish, DMA_start_address, 
      DMA_offset, DMA_read_write_filter_bias, DMA_filter_number, 
      \DMA_CNN_output_data[0][0] , \DMA_CNN_output_data[0][1] , 
      \DMA_CNN_output_data[0][2] , \DMA_CNN_output_data[0][3] , 
      \DMA_CNN_output_data[0][4] , \DMA_CNN_output_data[1][0] , 
      \DMA_CNN_output_data[1][1] , \DMA_CNN_output_data[1][2] , 
      \DMA_CNN_output_data[1][3] , \DMA_CNN_output_data[1][4] , 
      \DMA_CNN_output_data[2][0] , \DMA_CNN_output_data[2][1] , 
      \DMA_CNN_output_data[2][2] , \DMA_CNN_output_data[2][3] , 
      \DMA_CNN_output_data[2][4] , \DMA_CNN_output_data[3][0] , 
      \DMA_CNN_output_data[3][1] , \DMA_CNN_output_data[3][2] , 
      \DMA_CNN_output_data[3][3] , \DMA_CNN_output_data[3][4] , 
      \DMA_CNN_output_data[4][0] , \DMA_CNN_output_data[4][1] , 
      \DMA_CNN_output_data[4][2] , \DMA_CNN_output_data[4][3] , 
      \DMA_CNN_output_data[4][4] , DMA_CNN_input_data);
   input start;
   input reset;
   output finish;
   input clk;
   input [15:0]\filter[0][0] ;
   input [15:0]\filter[0][1] ;
   input [15:0]\filter[0][2] ;
   input [15:0]\filter[0][3] ;
   input [15:0]\filter[0][4] ;
   input [15:0]\filter[1][0] ;
   input [15:0]\filter[1][1] ;
   input [15:0]\filter[1][2] ;
   input [15:0]\filter[1][3] ;
   input [15:0]\filter[1][4] ;
   input [15:0]\filter[2][0] ;
   input [15:0]\filter[2][1] ;
   input [15:0]\filter[2][2] ;
   input [15:0]\filter[2][3] ;
   input [15:0]\filter[2][4] ;
   input [15:0]\filter[3][0] ;
   input [15:0]\filter[3][1] ;
   input [15:0]\filter[3][2] ;
   input [15:0]\filter[3][3] ;
   input [15:0]\filter[3][4] ;
   input [15:0]\filter[4][0] ;
   input [15:0]\filter[4][1] ;
   input [15:0]\filter[4][2] ;
   input [15:0]\filter[4][3] ;
   input [15:0]\filter[4][4] ;
   output [15:0]FB_index_bias;
   input [15:0]FB_output_bias;
   output [15:0]index_filter;
   output DMA_start;
   input DMA_finish;
   output [15:0]DMA_start_address;
   output [15:0]DMA_offset;
   output [1:0]DMA_read_write_filter_bias;
   output [15:0]DMA_filter_number;
   input [15:0]\DMA_CNN_output_data[0][0] ;
   input [15:0]\DMA_CNN_output_data[0][1] ;
   input [15:0]\DMA_CNN_output_data[0][2] ;
   input [15:0]\DMA_CNN_output_data[0][3] ;
   input [15:0]\DMA_CNN_output_data[0][4] ;
   input [15:0]\DMA_CNN_output_data[1][0] ;
   input [15:0]\DMA_CNN_output_data[1][1] ;
   input [15:0]\DMA_CNN_output_data[1][2] ;
   input [15:0]\DMA_CNN_output_data[1][3] ;
   input [15:0]\DMA_CNN_output_data[1][4] ;
   input [15:0]\DMA_CNN_output_data[2][0] ;
   input [15:0]\DMA_CNN_output_data[2][1] ;
   input [15:0]\DMA_CNN_output_data[2][2] ;
   input [15:0]\DMA_CNN_output_data[2][3] ;
   input [15:0]\DMA_CNN_output_data[2][4] ;
   input [15:0]\DMA_CNN_output_data[3][0] ;
   input [15:0]\DMA_CNN_output_data[3][1] ;
   input [15:0]\DMA_CNN_output_data[3][2] ;
   input [15:0]\DMA_CNN_output_data[3][3] ;
   input [15:0]\DMA_CNN_output_data[3][4] ;
   input [15:0]\DMA_CNN_output_data[4][0] ;
   input [15:0]\DMA_CNN_output_data[4][1] ;
   input [15:0]\DMA_CNN_output_data[4][2] ;
   input [15:0]\DMA_CNN_output_data[4][3] ;
   input [15:0]\DMA_CNN_output_data[4][4] ;
   output [15:0]DMA_CNN_input_data;

   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_230;
   wire n_0_231;
   wire n_0_232;
   wire n_0_233;
   wire n_0_235;
   wire n_0_236;
   wire n_0_237;
   wire n_0_238;
   wire n_0_239;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_248;
   wire n_0_249;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_256;
   wire n_0_257;
   wire n_0_258;
   wire n_0_259;
   wire n_0_260;
   wire n_0_261;
   wire n_0_295;
   wire n_0_296;
   wire n_0_297;
   wire n_0_298;
   wire n_0_299;
   wire n_0_300;
   wire n_0_301;
   wire n_0_302;
   wire n_0_303;
   wire n_0_304;
   wire n_0_305;
   wire n_0_306;
   wire n_0_307;
   wire n_0_308;
   wire n_0_309;
   wire n_0_310;
   wire n_0_311;
   wire n_0_312;
   wire n_0_313;
   wire n_0_314;
   wire n_0_315;
   wire n_0_316;
   wire n_0_317;
   wire n_0_318;
   wire n_0_319;
   wire n_0_320;
   wire n_0_321;
   wire n_0_322;
   wire n_0_323;
   wire n_0_324;
   wire n_0_325;
   wire n_0_326;
   wire n_0_327;
   wire n_0_328;
   wire n_0_329;
   wire n_0_330;
   wire n_0_331;
   wire n_0_332;
   wire n_0_333;
   wire n_0_334;
   wire n_0_335;
   wire n_0_336;
   wire n_0_337;
   wire n_0_338;
   wire n_0_339;
   wire n_0_340;
   wire n_0_341;
   wire n_0_342;
   wire n_0_343;
   wire n_0_363;
   wire n_0_364;
   wire n_0_365;
   wire n_0_366;
   wire n_0_367;
   wire n_0_368;
   wire n_0_369;
   wire n_0_370;
   wire n_0_371;
   wire n_0_372;
   wire n_0_373;
   wire n_0_374;
   wire n_0_375;
   wire n_0_376;
   wire n_0_377;
   wire n_0_378;
   wire n_0_379;
   wire n_0_380;
   wire n_0_381;
   wire n_0_382;
   wire n_0_383;
   wire n_0_384;
   wire n_0_385;
   wire n_0_386;
   wire n_0_387;
   wire n_0_388;
   wire n_0_389;
   wire n_0_390;
   wire n_0_391;
   wire n_0_392;
   wire n_0_393;
   wire n_0_394;
   wire n_0_395;
   wire n_0_396;
   wire n_0_397;
   wire n_0_398;
   wire n_0_399;
   wire n_0_400;
   wire n_0_401;
   wire n_0_402;
   wire n_0_403;
   wire n_0_404;
   wire n_0_405;
   wire n_0_406;
   wire n_0_407;
   wire n_0_408;
   wire n_0_409;
   wire n_0_410;
   wire n_0_411;
   wire n_0_412;
   wire n_0_413;
   wire n_0_414;
   wire n_0_415;
   wire n_0_416;
   wire n_0_417;
   wire n_0_418;
   wire n_0_419;
   wire n_0_420;
   wire n_0_421;
   wire n_0_422;
   wire n_0_423;
   wire n_0_424;
   wire n_0_425;
   wire n_0_426;
   wire n_0_427;
   wire n_0_428;
   wire n_0_429;
   wire n_0_430;
   wire n_0_431;
   wire n_0_432;
   wire n_0_433;
   wire n_0_434;
   wire n_0_435;
   wire n_0_436;
   wire n_0_437;
   wire n_0_438;
   wire n_0_440;
   wire n_0_441;
   wire n_0_458;
   wire n_0_459;
   wire n_0_460;
   wire n_0_461;
   wire n_0_462;
   wire n_0_463;
   wire n_0_464;
   wire n_0_465;
   wire n_0_466;
   wire n_0_467;
   wire n_0_468;
   wire n_0_469;
   wire n_0_470;
   wire n_0_471;
   wire n_0_472;
   wire n_0_473;
   wire n_0_474;
   wire n_0_475;
   wire n_0_476;
   wire n_0_477;
   wire n_0_478;
   wire n_0_479;
   wire n_0_480;
   wire n_0_481;
   wire n_0_482;
   wire n_0_483;
   wire n_0_484;
   wire n_0_485;
   wire n_0_486;
   wire n_0_2;
   wire [31:0]poolingState;
   wire [31:0]convResetState;
   wire convState;
   wire poolingReset;
   wire n_0_5;
   wire [31:0]layerCounter;
   wire writeReset;
   wire n_0_6;
   wire [15:0]writeAdress;
   wire n_0_7;
   wire [15:0]readAdress;
   wire convReset;
   wire n_0_8;
   wire [15:0]baseReadAdress;
   wire n_0_9;
   wire [31:0]kernelCounter;
   wire [31:0]filterCounter;
   wire n_0_14;
   wire [31:0]convWindowX;
   wire n_0_15;
   wire [31:0]poolingCounter;
   wire n_0_16;
   wire [31:0]poolingWindowX;
   wire n_0_510;
   wire [31:0]poolingWindowY;
   wire n_0_23;
   wire n_0_0_1;
   wire n_0_0_31;
   wire n_0_0_0;
   wire n_0_0_32;
   wire n_0_0_2;
   wire n_0_0_33;
   wire n_0_0_3;
   wire n_0_0_34;
   wire n_0_0_4;
   wire n_0_0_35;
   wire n_0_0_5;
   wire n_0_0_36;
   wire n_0_0_6;
   wire n_0_0_37;
   wire n_0_0_7;
   wire n_0_0_38;
   wire n_0_0_8;
   wire n_0_0_39;
   wire n_0_0_9;
   wire n_0_0_40;
   wire n_0_0_10;
   wire n_0_0_41;
   wire n_0_0_11;
   wire n_0_0_42;
   wire n_0_0_12;
   wire n_0_0_43;
   wire n_0_0_13;
   wire n_0_639;
   wire n_0_0_59;
   wire n_0_640;
   wire n_0_0_60;
   wire n_0_641;
   wire n_0_642;
   wire n_0_0_44;
   wire n_0_0_14;
   wire n_0_0_45;
   wire n_0_0_15;
   wire n_0_0_46;
   wire n_0_0_16;
   wire n_0_0_47;
   wire n_0_0_17;
   wire n_0_0_48;
   wire n_0_0_18;
   wire n_0_0_49;
   wire n_0_0_19;
   wire n_0_0_50;
   wire n_0_0_20;
   wire n_0_0_51;
   wire n_0_0_21;
   wire n_0_0_52;
   wire n_0_0_22;
   wire n_0_0_53;
   wire n_0_0_23;
   wire n_0_0_54;
   wire n_0_0_24;
   wire n_0_0_63;
   wire n_0_0_25;
   wire n_0_0_64;
   wire n_0_0_26;
   wire n_0_550;
   wire n_0_0_75;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_0_77;
   wire n_0_33;
   wire n_0_35;
   wire n_0_37;
   wire n_0_56;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_110;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_0_78;
   wire n_0_199;
   wire n_0_213;
   wire n_0_214;
   wire n_0_215;
   wire n_0_216;
   wire n_0_217;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_234;
   wire n_0_262;
   wire n_0_263;
   wire n_0_264;
   wire n_0_265;
   wire n_0_266;
   wire n_0_267;
   wire n_0_268;
   wire n_0_269;
   wire n_0_270;
   wire n_0_271;
   wire n_0_272;
   wire n_0_273;
   wire n_0_274;
   wire n_0_0_79;
   wire n_0_275;
   wire n_0_551;
   wire n_0_552;
   wire n_0_0_80;
   wire n_0_279;
   wire n_0_554;
   wire n_0_0_81;
   wire n_0_555;
   wire n_0_556;
   wire n_0_0_82;
   wire n_0_283;
   wire n_0_284;
   wire n_0_285;
   wire n_0_286;
   wire n_0_287;
   wire n_0_288;
   wire n_0_289;
   wire n_0_290;
   wire n_0_291;
   wire n_0_292;
   wire n_0_293;
   wire n_0_294;
   wire n_0_344;
   wire n_0_345;
   wire n_0_346;
   wire n_0_347;
   wire n_0_348;
   wire n_0_349;
   wire n_0_350;
   wire n_0_351;
   wire n_0_352;
   wire n_0_353;
   wire n_0_354;
   wire n_0_355;
   wire n_0_356;
   wire n_0_357;
   wire n_0_358;
   wire n_0_359;
   wire n_0_360;
   wire n_0_361;
   wire n_0_362;
   wire n_0_439;
   wire n_0_442;
   wire n_0_443;
   wire n_0_444;
   wire n_0_445;
   wire n_0_446;
   wire n_0_447;
   wire n_0_448;
   wire n_0_449;
   wire n_0_450;
   wire n_0_451;
   wire n_0_452;
   wire n_0_453;
   wire n_0_454;
   wire n_0_455;
   wire n_0_456;
   wire n_0_457;
   wire n_0_487;
   wire n_0_488;
   wire n_0_489;
   wire n_0_490;
   wire n_0_491;
   wire n_0_492;
   wire n_0_493;
   wire n_0_494;
   wire n_0_495;
   wire n_0_496;
   wire n_0_497;
   wire n_0_498;
   wire n_0_499;
   wire n_0_500;
   wire n_0_501;
   wire n_0_502;
   wire n_0_503;
   wire n_0_504;
   wire n_0_0;
   wire n_0_4;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_24;
   wire n_0_505;
   wire n_0_506;
   wire n_0_507;
   wire n_0_508;
   wire n_0_509;
   wire n_0_511;
   wire n_0_512;
   wire n_0_513;
   wire n_0_514;
   wire n_0_515;
   wire n_0_516;
   wire n_0_517;
   wire n_0_518;
   wire n_0_519;
   wire n_0_520;
   wire n_0_521;
   wire n_0_522;
   wire n_0_523;
   wire n_0_524;
   wire n_0_0_83;
   wire n_0_557;
   wire n_0_0_84;
   wire n_0_559;
   wire n_0_553;
   wire n_0_560;
   wire n_0_36;
   wire n_0_0_87;
   wire n_0_558;
   wire n_0_0_88;
   wire n_0_38;
   wire n_0_0_89;
   wire n_0_39;
   wire n_0_0_90;
   wire n_0_0_91;
   wire n_0_0_92;
   wire n_0_0_93;
   wire n_0_40;
   wire n_0_0_94;
   wire n_0_0_95;
   wire n_0_0_96;
   wire n_0_0_97;
   wire n_0_41;
   wire n_0_0_98;
   wire n_0_0_99;
   wire n_0_0_100;
   wire n_0_42;
   wire n_0_0_101;
   wire n_0_0_102;
   wire n_0_0_103;
   wire n_0_0_104;
   wire n_0_43;
   wire n_0_0_105;
   wire n_0_0_106;
   wire n_0_44;
   wire n_0_0_107;
   wire n_0_0_108;
   wire n_0_0_109;
   wire n_0_0_110;
   wire n_0_45;
   wire n_0_0_111;
   wire n_0_0_112;
   wire n_0_0_113;
   wire n_0_0_114;
   wire n_0_46;
   wire n_0_0_115;
   wire n_0_0_116;
   wire n_0_0_117;
   wire n_0_47;
   wire n_0_0_118;
   wire n_0_48;
   wire n_0_0_119;
   wire n_0_0_120;
   wire n_0_49;
   wire n_0_0_121;
   wire n_0_0_122;
   wire n_0_0_123;
   wire n_0_50;
   wire n_0_0_124;
   wire n_0_51;
   wire n_0_0_125;
   wire n_0_52;
   wire n_0_0_126;
   wire n_0_0_127;
   wire n_0_0_128;
   wire n_0_53;
   wire n_0_0_129;
   wire n_0_0_130;
   wire n_0_0_131;
   wire n_0_0_132;
   wire n_0_0_133;
   wire n_0_0_134;
   wire n_0_0_135;
   wire n_0_561;
   wire n_0_562;
   wire n_0_0_136;
   wire n_0_54;
   wire n_0_0_137;
   wire n_0_0_138;
   wire n_0_55;
   wire n_0_0_139;
   wire n_0_0_140;
   wire n_0_0_141;
   wire n_0_276;
   wire n_0_0_142;
   wire n_0_0_143;
   wire n_0_277;
   wire n_0_0_144;
   wire n_0_0_145;
   wire n_0_278;
   wire n_0_0_146;
   wire n_0_0_147;
   wire n_0_280;
   wire n_0_0_148;
   wire n_0_0_149;
   wire n_0_281;
   wire n_0_0_150;
   wire n_0_0_151;
   wire n_0_282;
   wire n_0_0_152;
   wire n_0_0_153;
   wire n_0_525;
   wire n_0_0_154;
   wire n_0_0_155;
   wire n_0_526;
   wire n_0_0_156;
   wire n_0_0_157;
   wire n_0_527;
   wire n_0_0_158;
   wire n_0_0_159;
   wire n_0_528;
   wire n_0_0_160;
   wire n_0_0_161;
   wire n_0_529;
   wire n_0_0_162;
   wire n_0_0_163;
   wire n_0_530;
   wire n_0_0_164;
   wire n_0_0_165;
   wire n_0_531;
   wire n_0_0_166;
   wire n_0_0_167;
   wire n_0_532;
   wire n_0_0_168;
   wire n_0_0_169;
   wire n_0_0_170;
   wire n_0_0_171;
   wire n_0_0_172;
   wire n_0_0_173;
   wire n_0_0_174;
   wire n_0_0_175;
   wire n_0_0_176;
   wire n_0_0_177;
   wire n_0_0_178;
   wire n_0_0_179;
   wire n_0_697;
   wire n_0_0_180;
   wire n_0_698;
   wire n_0_0_181;
   wire n_0_699;
   wire n_0_0_182;
   wire n_0_1;
   wire n_0_3;
   wire n_0_25;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_34;
   wire n_0_533;
   wire n_0_534;
   wire n_0_535;
   wire n_0_536;
   wire n_0_537;
   wire n_0_538;
   wire n_0_0_183;
   wire n_0_0_184;
   wire n_0_665;
   wire n_0_666;
   wire n_0_0_185;
   wire n_0_0_186;
   wire n_0_667;
   wire n_0_0_187;
   wire n_0_668;
   wire n_0_0_188;
   wire n_0_0_189;
   wire n_0_669;
   wire n_0_0_190;
   wire n_0_670;
   wire n_0_0_191;
   wire n_0_671;
   wire n_0_0_192;
   wire n_0_672;
   wire n_0_0_193;
   wire n_0_673;
   wire n_0_0_194;
   wire n_0_674;
   wire n_0_0_195;
   wire n_0_675;
   wire n_0_0_196;
   wire n_0_676;
   wire n_0_0_197;
   wire n_0_677;
   wire n_0_0_198;
   wire n_0_678;
   wire n_0_0_199;
   wire n_0_0_200;
   wire n_0_679;
   wire n_0_0_201;
   wire n_0_680;
   wire n_0_0_202;
   wire n_0_0_203;
   wire n_0_0_204;
   wire n_0_649;
   wire n_0_650;
   wire n_0_651;
   wire n_0_652;
   wire n_0_653;
   wire n_0_654;
   wire n_0_655;
   wire n_0_656;
   wire n_0_657;
   wire n_0_0_205;
   wire n_0_658;
   wire n_0_659;
   wire n_0_660;
   wire n_0_0_206;
   wire n_0_661;
   wire n_0_0_207;
   wire n_0_662;
   wire n_0_663;
   wire n_0_664;
   wire n_0_638;
   wire n_0_0_208;
   wire n_0_564;
   wire n_0_0_209;
   wire n_0_563;
   wire n_0_0_210;
   wire n_0_635;
   wire n_0_0_211;
   wire n_0_565;
   wire n_0_566;
   wire n_0_0_212;
   wire n_0_0_213;
   wire n_0_0_214;
   wire n_0_0_215;
   wire n_0_617;
   wire n_0_0_216;
   wire n_0_0_217;
   wire n_0_618;
   wire n_0_0_218;
   wire n_0_619;
   wire n_0_0_219;
   wire n_0_0_220;
   wire n_0_620;
   wire n_0_0_221;
   wire n_0_621;
   wire n_0_0_222;
   wire n_0_622;
   wire n_0_0_223;
   wire n_0_623;
   wire n_0_0_224;
   wire n_0_624;
   wire n_0_0_225;
   wire n_0_0_226;
   wire n_0_625;
   wire n_0_0_227;
   wire n_0_626;
   wire n_0_0_228;
   wire n_0_627;
   wire n_0_0_229;
   wire n_0_0_230;
   wire n_0_628;
   wire n_0_0_231;
   wire n_0_629;
   wire n_0_0_232;
   wire n_0_630;
   wire n_0_0_233;
   wire n_0_631;
   wire n_0_0_234;
   wire n_0_632;
   wire n_0_0_235;
   wire n_0_0_236;
   wire n_0_0_237;
   wire n_0_0_238;
   wire n_0_0_239;
   wire n_0_0_240;
   wire n_0_0_241;
   wire n_0_0_242;
   wire n_0_0_243;
   wire n_0_0_244;
   wire n_0_0_245;
   wire n_0_601;
   wire n_0_602;
   wire n_0_603;
   wire n_0_604;
   wire n_0_605;
   wire n_0_606;
   wire n_0_607;
   wire n_0_608;
   wire n_0_609;
   wire n_0_610;
   wire n_0_611;
   wire n_0_612;
   wire n_0_613;
   wire n_0_614;
   wire n_0_0_246;
   wire n_0_615;
   wire n_0_616;
   wire n_0_585;
   wire n_0_0_247;
   wire n_0_586;
   wire n_0_0_248;
   wire n_0_587;
   wire n_0_588;
   wire n_0_589;
   wire n_0_0_249;
   wire n_0_590;
   wire n_0_0_250;
   wire n_0_591;
   wire n_0_592;
   wire n_0_0_251;
   wire n_0_593;
   wire n_0_0_252;
   wire n_0_594;
   wire n_0_0_253;
   wire n_0_595;
   wire n_0_0_254;
   wire n_0_0_255;
   wire n_0_0_256;
   wire n_0_596;
   wire n_0_597;
   wire n_0_598;
   wire n_0_599;
   wire n_0_0_257;
   wire n_0_600;
   wire n_0_0_258;
   wire n_0_584;
   wire n_0_0_260;
   wire n_0_0_261;
   wire n_0_0_262;
   wire n_0_0_263;
   wire n_0_0_264;
   wire n_0_0_265;
   wire n_0_0_266;
   wire n_0_0_267;
   wire n_0_0_268;
   wire n_0_567;
   wire n_0_0_269;
   wire n_0_0_270;
   wire n_0_0_271;
   wire n_0_0_272;
   wire n_0_0_273;
   wire n_0_0_274;
   wire n_0_0_275;
   wire n_0_0_276;
   wire n_0_0_277;
   wire n_0_0_278;
   wire n_0_568;
   wire n_0_569;
   wire n_0_0_280;
   wire n_0_0_281;
   wire n_0_0_282;
   wire n_0_0_283;
   wire n_0_0_284;
   wire n_0_0_285;
   wire n_0_0_286;
   wire n_0_0_287;
   wire n_0_0_288;
   wire n_0_0_289;
   wire n_0_0_290;
   wire n_0_0_291;
   wire n_0_0_292;
   wire n_0_0_293;
   wire n_0_0_294;
   wire n_0_0_295;
   wire n_0_0_296;
   wire n_0_0_297;
   wire n_0_0_298;
   wire n_0_0_299;
   wire n_0_0_300;
   wire n_0_0_301;
   wire n_0_0_302;
   wire n_0_0_303;
   wire n_0_0_304;
   wire n_0_0_305;
   wire n_0_0_306;
   wire n_0_0_307;
   wire n_0_0_308;
   wire n_0_0_309;
   wire n_0_0_310;
   wire n_0_0_311;
   wire n_0_0_312;
   wire n_0_0_313;
   wire n_0_0_314;
   wire n_0_0_315;
   wire n_0_0_316;
   wire n_0_0_317;
   wire n_0_0_318;
   wire n_0_0_319;
   wire n_0_0_320;
   wire n_0_0_321;
   wire n_0_0_322;
   wire n_0_0_323;
   wire n_0_0_324;
   wire n_0_0_325;
   wire n_0_0_326;
   wire n_0_0_327;
   wire n_0_0_328;
   wire n_0_0_329;
   wire n_0_0_330;
   wire n_0_0_331;
   wire n_0_0_332;
   wire n_0_0_333;
   wire n_0_0_334;
   wire n_0_0_335;
   wire n_0_0_336;
   wire n_0_0_337;
   wire n_0_0_338;
   wire n_0_0_339;
   wire n_0_0_340;
   wire n_0_0_341;
   wire n_0_0_342;
   wire n_0_0_343;
   wire n_0_0_344;
   wire n_0_0_345;
   wire n_0_0_346;
   wire n_0_0_347;
   wire n_0_0_348;
   wire n_0_0_349;
   wire n_0_0_350;
   wire n_0_0_351;
   wire n_0_0_352;
   wire n_0_0_353;
   wire n_0_0_354;
   wire n_0_0_355;
   wire n_0_0_356;
   wire n_0_0_357;
   wire n_0_0_358;
   wire n_0_0_359;
   wire n_0_0_360;
   wire n_0_0_361;
   wire n_0_0_362;
   wire n_0_0_363;
   wire n_0_0_364;
   wire n_0_0_365;
   wire n_0_0_366;
   wire n_0_0_367;
   wire n_0_0_368;
   wire n_0_0_369;
   wire n_0_0_370;
   wire n_0_0_371;
   wire n_0_0_372;
   wire n_0_0_373;
   wire n_0_0_374;
   wire n_0_0_375;
   wire n_0_0_376;
   wire n_0_0_377;
   wire n_0_0_378;
   wire n_0_0_379;
   wire n_0_0_380;
   wire n_0_0_381;
   wire n_0_0_382;
   wire n_0_0_383;
   wire n_0_0_384;
   wire n_0_0_385;
   wire n_0_0_386;
   wire n_0_0_387;
   wire n_0_0_388;
   wire n_0_0_389;
   wire n_0_0_390;
   wire n_0_0_391;
   wire n_0_0_392;
   wire n_0_0_394;
   wire n_0_0_398;
   wire n_0_0_399;
   wire n_0_0_400;
   wire n_0_0_401;
   wire n_0_0_402;
   wire n_0_0_403;
   wire n_0_0_404;
   wire n_0_0_405;
   wire n_0_0_406;
   wire n_0_0_407;
   wire n_0_0_408;
   wire n_0_0_409;
   wire n_0_0_410;
   wire n_0_0_411;
   wire n_0_0_412;
   wire n_0_0_413;
   wire n_0_0_414;
   wire n_0_0_415;
   wire n_0_0_416;
   wire n_0_0_417;
   wire n_0_0_418;
   wire n_0_0_419;
   wire n_0_0_420;
   wire n_0_0_421;
   wire n_0_0_422;
   wire n_0_0_423;
   wire n_0_0_424;
   wire n_0_0_425;
   wire n_0_0_426;
   wire n_0_0_427;
   wire n_0_573;
   wire n_0_0_428;
   wire n_0_0_430;
   wire n_0_0_431;
   wire n_0_0_432;
   wire n_0_0_433;
   wire n_0_549;
   wire n_0_0_434;
   wire n_0_0_435;
   wire n_0_540;
   wire n_0_539;
   wire n_0_541;
   wire n_0_0_436;
   wire n_0_542;
   wire n_0_0_437;
   wire n_0_543;
   wire n_0_544;
   wire n_0_545;
   wire n_0_546;
   wire n_0_547;
   wire n_0_0_27;
   wire n_0_0_438;
   wire n_0_0_439;
   wire n_0_0_440;
   wire n_0_0_441;
   wire n_0_570;
   wire n_0_0_442;
   wire n_0_681;
   wire n_0_682;
   wire n_0_683;
   wire n_0_684;
   wire n_0_685;
   wire n_0_0_28;
   wire n_0_686;
   wire n_0_0_29;
   wire n_0_687;
   wire n_0_0_30;
   wire n_0_688;
   wire n_0_0_55;
   wire n_0_689;
   wire n_0_0_443;
   wire n_0_690;
   wire n_0_0_56;
   wire n_0_691;
   wire n_0_0_57;
   wire n_0_692;
   wire n_0_0_58;
   wire n_0_0_444;
   wire n_0_0_445;
   wire n_0_0_446;
   wire n_0_693;
   wire n_0_0_447;
   wire n_0_694;
   wire n_0_0_61;
   wire n_0_0_448;
   wire n_0_0_449;
   wire n_0_0_450;
   wire n_0_0_451;
   wire n_0_695;
   wire n_0_696;
   wire n_0_644;
   wire n_0_0_452;
   wire n_0_645;
   wire n_0_583;
   wire n_0_581;
   wire n_0_0_453;
   wire n_0_0_454;
   wire n_0_571;
   wire n_0_0_455;
   wire n_0_548;
   wire n_0_0_456;
   wire n_0_0_62;
   wire n_0_0_457;
   wire n_0_0_458;
   wire n_0_0_459;
   wire n_0_0_460;
   wire n_0_0_461;
   wire n_0_572;
   wire n_0_0_462;
   wire n_0_646;
   wire n_0_0_463;
   wire n_0_0_65;
   wire n_0_0_464;
   wire n_0_0_465;
   wire n_0_0_466;
   wire n_0_0_467;
   wire n_0_0_468;
   wire n_0_0_469;
   wire n_0_0_470;
   wire n_0_0_471;
   wire n_0_0_472;
   wire n_0_0_473;
   wire n_0_0_474;
   wire n_0_0_475;
   wire n_0_0_66;
   wire n_0_0_67;
   wire n_0_0_68;
   wire n_0_0_69;
   wire n_0_0_70;
   wire n_0_0_71;
   wire n_0_0_72;
   wire n_0_0_73;
   wire n_0_0_74;
   wire n_0_0_76;
   wire n_0_0_85;
   wire n_0_0_86;
   wire n_0_0_259;
   wire n_0_0_279;
   wire n_0_0_393;
   wire n_0_0_395;
   wire n_0_0_396;
   wire n_0_0_397;
   wire n_0_0_429;
   wire n_0_576;
   wire n_0_575;
   wire n_0_574;
   wire n_0_578;
   wire n_0_577;
   wire n_0_579;
   wire n_0_580;
   wire n_0_633;
   wire n_0_582;
   wire n_0_636;
   wire n_0_634;
   wire n_0_637;
   wire n_0_643;
   wire n_0_647;
   wire n_0_648;

   datapath__0_4270 i_0_36 (.p_0({n_0_600, n_0_599, n_0_598, n_0_597, n_0_596, 
      n_0_595, n_0_594, n_0_593, n_0_592, n_0_591, n_0_590, n_0_589, n_0_588, 
      n_0_587, n_0_586, n_0_585}), .p_1({n_0_71, n_0_70, n_0_69, n_0_68, n_0_67, 
      n_0_66, n_0_65, n_0_64, n_0_63, n_0_62, n_0_61, n_0_60, n_0_59, n_0_58, 
      n_0_57, uc_0}));
   datapath__0_4273 i_0_39 (.p_0({n_0_616, n_0_615, n_0_614, n_0_613, n_0_612, 
      n_0_611, n_0_610, n_0_609, n_0_608, n_0_607, n_0_606, n_0_605, n_0_604, 
      n_0_603, n_0_602, n_0_601}), .p_1({n_0_93, n_0_92, n_0_91, n_0_90, n_0_89, 
      n_0_88, n_0_87, n_0_86, n_0_85, n_0_84, n_0_83, n_0_82, n_0_81, n_0_80, 
      n_0_79, n_0_78}));
   datapath__0_4284 i_0_50 (.p_0({n_0_664, n_0_663, n_0_662, n_0_661, n_0_660, 
      n_0_659, n_0_658, n_0_657, n_0_656, n_0_655, n_0_654, n_0_653, n_0_652, 
      n_0_651, n_0_650, n_0_649}), .p_1({n_0_109, n_0_108, n_0_107, n_0_106, 
      n_0_105, n_0_104, n_0_103, n_0_102, n_0_101, n_0_100, n_0_99, n_0_98, 
      n_0_97, n_0_96, n_0_95, n_0_94}));
   datapath__0_4288 i_0_53 (.featureMapSize({1'b0, n_0_570, n_0_581, n_0_646, 
      n_0_645, n_0_548, n_0_644}), .p_0({n_0_696, n_0_695, n_0_694, n_0_693, 
      n_0_692, n_0_691, n_0_690, n_0_689, n_0_688, n_0_687, n_0_686, n_0_685, 
      n_0_684, n_0_683, n_0_682, n_0_681}), .p_1({n_0_136, n_0_135, n_0_134, 
      n_0_133, n_0_132, n_0_131, n_0_130, n_0_119, n_0_118, n_0_117, n_0_116, 
      n_0_115, n_0_114, n_0_113, n_0_112, n_0_111}));
   datapath__0_4294 i_0_59 (.p_0({n_0_547, n_0_546, n_0_545, n_0_544, n_0_543, 
      n_0_542, n_0_541, n_0_540, n_0_539, uc_1, n_0_644}), .p_1({n_0_109, 
      n_0_108, n_0_107, n_0_106, n_0_105, n_0_104, n_0_103, n_0_102, n_0_101, 
      n_0_100, n_0_99, n_0_98, n_0_97, n_0_96, n_0_95, n_0_94}), .p_2({n_0_180, 
      n_0_179, n_0_178, n_0_177, n_0_176, n_0_175, n_0_174, n_0_173, n_0_172, 
      n_0_171, n_0_170, n_0_169, n_0_168, n_0_167, n_0_166, n_0_165}));
   datapath__0_4295 i_0_60 (.p_0({uc_2, n_0_570, n_0_581, n_0_642, n_0_641, 
      n_0_640, n_0_639, n_0_583, n_0_572, n_0_548, 1'b0, n_0_644}), .p_1({
      n_0_538, n_0_537, n_0_536, n_0_535, n_0_534, n_0_533, n_0_34, n_0_32, 
      n_0_31, n_0_30, n_0_25, n_0_3, n_0_1, n_0_699, n_0_698, n_0_697}), 
      .p_2({n_0_212, n_0_211, n_0_210, n_0_209, n_0_208, n_0_207, n_0_206, 
      n_0_205, n_0_204, n_0_203, n_0_202, n_0_201, n_0_200, n_0_183, n_0_182, 
      n_0_181}));
   datapath__0_4312 i_0_77 (.filterCounter(filterCounter), .p_0({n_0_261, 
      n_0_260, n_0_259, n_0_258, n_0_257, n_0_256, n_0_255, n_0_254, n_0_253, 
      n_0_252, n_0_251, n_0_250, n_0_249, n_0_248, n_0_247, n_0_246, n_0_245, 
      n_0_244, n_0_243, n_0_242, n_0_241, n_0_240, n_0_239, n_0_238, n_0_237, 
      n_0_236, n_0_235, n_0_233, n_0_232, n_0_231, n_0_230, uc_3}));
   datapath__0_4318 i_0_83 (.convWindowX(convWindowX), .p_0({n_0_325, n_0_324, 
      n_0_323, n_0_322, n_0_321, n_0_320, n_0_319, n_0_318, n_0_317, n_0_316, 
      n_0_315, n_0_314, n_0_313, n_0_312, n_0_311, n_0_310, n_0_309, n_0_308, 
      n_0_307, n_0_306, n_0_305, n_0_304, n_0_303, n_0_302, n_0_301, n_0_300, 
      n_0_299, n_0_298, n_0_297, n_0_296, n_0_295, uc_4}));
   datapath__0_4321 i_0_86 (.kernelCounter(kernelCounter), .p_0({n_0_376, 
      n_0_375, n_0_374, n_0_373, n_0_372, n_0_371, n_0_370, n_0_369, n_0_368, 
      n_0_367, n_0_366, n_0_365, n_0_364, n_0_363, n_0_343, n_0_342, n_0_341, 
      n_0_340, n_0_339, n_0_338, n_0_337, n_0_336, n_0_335, n_0_334, n_0_333, 
      n_0_332, n_0_331, n_0_330, n_0_329, n_0_328, n_0_327, n_0_326}));
   datapath__0_4332 i_0_97 (.poolingWindowY({poolingWindowY[31], 
      poolingWindowY[30], poolingWindowY[29], poolingWindowY[28], 
      poolingWindowY[27], poolingWindowY[26], poolingWindowY[25], 
      poolingWindowY[24], poolingWindowY[23], poolingWindowY[22], 
      poolingWindowY[21], poolingWindowY[20], poolingWindowY[19], 
      poolingWindowY[18], poolingWindowY[17], poolingWindowY[16], 
      poolingWindowY[15], poolingWindowY[14], poolingWindowY[13], 
      poolingWindowY[12], poolingWindowY[11], poolingWindowY[10], 
      poolingWindowY[9], poolingWindowY[8], poolingWindowY[7], poolingWindowY[6], 
      poolingWindowY[5], poolingWindowY[4], poolingWindowY[3], poolingWindowY[2], 
      poolingWindowY[1], uc_5}), .p_0({n_0_407, n_0_406, n_0_405, n_0_404, 
      n_0_403, n_0_402, n_0_401, n_0_400, n_0_399, n_0_398, n_0_397, n_0_396, 
      n_0_395, n_0_394, n_0_393, n_0_392, n_0_391, n_0_390, n_0_389, n_0_388, 
      n_0_387, n_0_386, n_0_385, n_0_384, n_0_383, n_0_382, n_0_381, n_0_380, 
      n_0_379, n_0_378, n_0_377, uc_6}));
   datapath__0_4335 i_0_100 (.poolingWindowX({poolingWindowX[31], 
      poolingWindowX[30], poolingWindowX[29], poolingWindowX[28], 
      poolingWindowX[27], poolingWindowX[26], poolingWindowX[25], 
      poolingWindowX[24], poolingWindowX[23], poolingWindowX[22], 
      poolingWindowX[21], poolingWindowX[20], poolingWindowX[19], 
      poolingWindowX[18], poolingWindowX[17], poolingWindowX[16], 
      poolingWindowX[15], poolingWindowX[14], poolingWindowX[13], 
      poolingWindowX[12], poolingWindowX[11], poolingWindowX[10], 
      poolingWindowX[9], poolingWindowX[8], poolingWindowX[7], poolingWindowX[6], 
      poolingWindowX[5], poolingWindowX[4], poolingWindowX[3], poolingWindowX[2], 
      poolingWindowX[1], uc_7}), .p_0({n_0_438, n_0_437, n_0_436, n_0_435, 
      n_0_434, n_0_433, n_0_432, n_0_431, n_0_430, n_0_429, n_0_428, n_0_427, 
      n_0_426, n_0_425, n_0_424, n_0_423, n_0_422, n_0_421, n_0_420, n_0_419, 
      n_0_418, n_0_417, n_0_416, n_0_415, n_0_414, n_0_413, n_0_412, n_0_411, 
      n_0_410, n_0_409, n_0_408, uc_8}));
   datapath__0_4338 i_0_103 (.poolingCounter(poolingCounter), .p_0({n_0_486, 
      n_0_485, n_0_484, n_0_483, n_0_482, n_0_481, n_0_480, n_0_479, n_0_478, 
      n_0_477, n_0_476, n_0_475, n_0_474, n_0_473, n_0_472, n_0_471, n_0_470, 
      n_0_469, n_0_468, n_0_467, n_0_466, n_0_465, n_0_464, n_0_463, n_0_462, 
      n_0_461, n_0_460, n_0_459, n_0_458, n_0_441, n_0_440, uc_9}));
   DFF_X1 \DMA_filter_number_reg[2]  (.D(n_0_576), .CK(clk), .Q(
      DMA_filter_number[2]), .QN());
   DFF_X1 \DMA_filter_number_reg[6]  (.D(n_0_575), .CK(clk), .Q(
      DMA_filter_number[6]), .QN());
   DFF_X1 \DMA_filter_number_reg[10]  (.D(n_0_574), .CK(clk), .Q(
      DMA_filter_number[10]), .QN());
   DFF_X1 \DMA_read_write_filter_bias_reg[0]  (.D(n_0_578), .CK(clk), .Q(
      DMA_read_write_filter_bias[0]), .QN());
   DFF_X1 \DMA_read_write_filter_bias_reg[1]  (.D(n_0_577), .CK(clk), .Q(
      DMA_read_write_filter_bias[1]), .QN());
   CLKGATETST_X1 clk_gate_DMA_start_address_reg (.CK(clk), .E(n_0_569), .SE(1'b0), 
      .GCK(n_0_2));
   DFF_X1 \DMA_start_address_reg[15]  (.D(n_0_53), .CK(n_0_2), .Q(
      DMA_start_address[15]), .QN());
   DFF_X1 \DMA_start_address_reg[14]  (.D(n_0_52), .CK(n_0_2), .Q(
      DMA_start_address[14]), .QN());
   DFF_X1 \DMA_start_address_reg[13]  (.D(n_0_51), .CK(n_0_2), .Q(
      DMA_start_address[13]), .QN());
   DFF_X1 \DMA_start_address_reg[12]  (.D(n_0_50), .CK(n_0_2), .Q(
      DMA_start_address[12]), .QN());
   DFF_X1 \DMA_start_address_reg[11]  (.D(n_0_49), .CK(n_0_2), .Q(
      DMA_start_address[11]), .QN());
   DFF_X1 \DMA_start_address_reg[10]  (.D(n_0_48), .CK(n_0_2), .Q(
      DMA_start_address[10]), .QN());
   DFF_X1 \DMA_start_address_reg[9]  (.D(n_0_47), .CK(n_0_2), .Q(
      DMA_start_address[9]), .QN());
   DFF_X1 \DMA_start_address_reg[8]  (.D(n_0_46), .CK(n_0_2), .Q(
      DMA_start_address[8]), .QN());
   DFF_X1 \DMA_start_address_reg[7]  (.D(n_0_45), .CK(n_0_2), .Q(
      DMA_start_address[7]), .QN());
   DFF_X1 \DMA_start_address_reg[6]  (.D(n_0_44), .CK(n_0_2), .Q(
      DMA_start_address[6]), .QN());
   DFF_X1 \DMA_start_address_reg[5]  (.D(n_0_43), .CK(n_0_2), .Q(
      DMA_start_address[5]), .QN());
   DFF_X1 \DMA_start_address_reg[4]  (.D(n_0_42), .CK(n_0_2), .Q(
      DMA_start_address[4]), .QN());
   DFF_X1 \DMA_start_address_reg[3]  (.D(n_0_41), .CK(n_0_2), .Q(
      DMA_start_address[3]), .QN());
   DFF_X1 \DMA_start_address_reg[2]  (.D(n_0_40), .CK(n_0_2), .Q(
      DMA_start_address[2]), .QN());
   DFF_X1 \DMA_start_address_reg[1]  (.D(n_0_39), .CK(n_0_2), .Q(
      DMA_start_address[1]), .QN());
   DFF_X1 \DMA_start_address_reg[0]  (.D(n_0_38), .CK(n_0_2), .Q(
      DMA_start_address[0]), .QN());
   DFF_X1 finishCNN_reg (.D(n_0_579), .CK(clk), .Q(finish), .QN());
   DFF_X1 DMA_start_reg (.D(n_0_580), .CK(clk), .Q(DMA_start), .QN());
   DFF_X1 \poolingState_reg[0]  (.D(n_0_633), .CK(clk), .Q(poolingState[0]), 
      .QN());
   DFF_X1 \poolingState_reg[1]  (.D(n_0_582), .CK(clk), .Q(poolingState[1]), 
      .QN());
   DFF_X1 \convResetState_reg[0]  (.D(n_0_636), .CK(clk), .Q(convResetState[0]), 
      .QN());
   DFF_X1 \convResetState_reg[1]  (.D(n_0_634), .CK(clk), .Q(convResetState[1]), 
      .QN());
   DFF_X1 convState_reg (.D(n_0_637), .CK(clk), .Q(convState), .QN());
   DFF_X1 poolingReset_reg (.D(n_0_643), .CK(clk), .Q(poolingReset), .QN());
   CLKGATETST_X1 clk_gate_layerCounter_reg (.CK(clk), .E(n_0_279), .SE(1'b0), 
      .GCK(n_0_5));
   DFF_X1 \layerCounter_reg[31]  (.D(n_0_29), .CK(n_0_5), .Q(layerCounter[31]), 
      .QN());
   DFF_X1 \layerCounter_reg[2]  (.D(n_0_28), .CK(n_0_5), .Q(layerCounter[2]), 
      .QN());
   DFF_X1 \layerCounter_reg[1]  (.D(n_0_27), .CK(n_0_5), .Q(layerCounter[1]), 
      .QN());
   DFF_X1 \layerCounter_reg[0]  (.D(n_0_26), .CK(n_0_5), .Q(layerCounter[0]), 
      .QN());
   DFF_X1 writeReset_reg (.D(n_0_647), .CK(clk), .Q(writeReset), .QN());
   CLKGATETST_X1 clk_gate_writeAdress_reg (.CK(clk), .E(n_0_584), .SE(1'b0), 
      .GCK(n_0_6));
   DFF_X1 \writeAdress_reg[15]  (.D(n_0_632), .CK(n_0_6), .Q(writeAdress[15]), 
      .QN());
   DFF_X1 \writeAdress_reg[14]  (.D(n_0_631), .CK(n_0_6), .Q(writeAdress[14]), 
      .QN());
   DFF_X1 \writeAdress_reg[13]  (.D(n_0_630), .CK(n_0_6), .Q(writeAdress[13]), 
      .QN());
   DFF_X1 \writeAdress_reg[12]  (.D(n_0_629), .CK(n_0_6), .Q(writeAdress[12]), 
      .QN());
   DFF_X1 \writeAdress_reg[11]  (.D(n_0_628), .CK(n_0_6), .Q(writeAdress[11]), 
      .QN());
   DFF_X1 \writeAdress_reg[10]  (.D(n_0_627), .CK(n_0_6), .Q(writeAdress[10]), 
      .QN());
   DFF_X1 \writeAdress_reg[9]  (.D(n_0_626), .CK(n_0_6), .Q(writeAdress[9]), 
      .QN());
   DFF_X1 \writeAdress_reg[8]  (.D(n_0_625), .CK(n_0_6), .Q(writeAdress[8]), 
      .QN());
   DFF_X1 \writeAdress_reg[7]  (.D(n_0_624), .CK(n_0_6), .Q(writeAdress[7]), 
      .QN());
   DFF_X1 \writeAdress_reg[6]  (.D(n_0_623), .CK(n_0_6), .Q(writeAdress[6]), 
      .QN());
   DFF_X1 \writeAdress_reg[5]  (.D(n_0_622), .CK(n_0_6), .Q(writeAdress[5]), 
      .QN());
   DFF_X1 \writeAdress_reg[4]  (.D(n_0_621), .CK(n_0_6), .Q(writeAdress[4]), 
      .QN());
   DFF_X1 \writeAdress_reg[3]  (.D(n_0_620), .CK(n_0_6), .Q(writeAdress[3]), 
      .QN());
   DFF_X1 \writeAdress_reg[2]  (.D(n_0_619), .CK(n_0_6), .Q(writeAdress[2]), 
      .QN());
   DFF_X1 \writeAdress_reg[1]  (.D(n_0_618), .CK(n_0_6), .Q(writeAdress[1]), 
      .QN());
   DFF_X1 \writeAdress_reg[0]  (.D(n_0_617), .CK(n_0_6), .Q(writeAdress[0]), 
      .QN());
   CLKGATETST_X1 clk_gate_readAdress_reg (.CK(clk), .E(n_0_635), .SE(1'b0), 
      .GCK(n_0_7));
   DFF_X1 \readAdress_reg[15]  (.D(n_0_532), .CK(n_0_7), .Q(readAdress[15]), 
      .QN());
   DFF_X1 \readAdress_reg[14]  (.D(n_0_531), .CK(n_0_7), .Q(readAdress[14]), 
      .QN());
   DFF_X1 \readAdress_reg[13]  (.D(n_0_530), .CK(n_0_7), .Q(readAdress[13]), 
      .QN());
   DFF_X1 \readAdress_reg[12]  (.D(n_0_529), .CK(n_0_7), .Q(readAdress[12]), 
      .QN());
   DFF_X1 \readAdress_reg[11]  (.D(n_0_528), .CK(n_0_7), .Q(readAdress[11]), 
      .QN());
   DFF_X1 \readAdress_reg[10]  (.D(n_0_527), .CK(n_0_7), .Q(readAdress[10]), 
      .QN());
   DFF_X1 \readAdress_reg[9]  (.D(n_0_526), .CK(n_0_7), .Q(readAdress[9]), .QN());
   DFF_X1 \readAdress_reg[8]  (.D(n_0_525), .CK(n_0_7), .Q(readAdress[8]), .QN());
   DFF_X1 \readAdress_reg[7]  (.D(n_0_282), .CK(n_0_7), .Q(readAdress[7]), .QN());
   DFF_X1 \readAdress_reg[6]  (.D(n_0_281), .CK(n_0_7), .Q(readAdress[6]), .QN());
   DFF_X1 \readAdress_reg[5]  (.D(n_0_280), .CK(n_0_7), .Q(readAdress[5]), .QN());
   DFF_X1 \readAdress_reg[4]  (.D(n_0_278), .CK(n_0_7), .Q(readAdress[4]), .QN());
   DFF_X1 \readAdress_reg[3]  (.D(n_0_277), .CK(n_0_7), .Q(readAdress[3]), .QN());
   DFF_X1 \readAdress_reg[2]  (.D(n_0_276), .CK(n_0_7), .Q(readAdress[2]), .QN());
   DFF_X1 \readAdress_reg[1]  (.D(n_0_55), .CK(n_0_7), .Q(readAdress[1]), .QN());
   DFF_X1 \readAdress_reg[0]  (.D(n_0_54), .CK(n_0_7), .Q(readAdress[0]), .QN());
   DFF_X1 convReset_reg (.D(n_0_648), .CK(clk), .Q(convReset), .QN());
   CLKGATETST_X1 clk_gate_baseReadAdress_reg (.CK(clk), .E(n_0_638), .SE(1'b0), 
      .GCK(n_0_8));
   DFF_X1 \baseReadAdress_reg[15]  (.D(n_0_680), .CK(n_0_8), .Q(
      baseReadAdress[15]), .QN());
   DFF_X1 \baseReadAdress_reg[14]  (.D(n_0_679), .CK(n_0_8), .Q(
      baseReadAdress[14]), .QN());
   DFF_X1 \baseReadAdress_reg[13]  (.D(n_0_678), .CK(n_0_8), .Q(
      baseReadAdress[13]), .QN());
   DFF_X1 \baseReadAdress_reg[12]  (.D(n_0_677), .CK(n_0_8), .Q(
      baseReadAdress[12]), .QN());
   DFF_X1 \baseReadAdress_reg[11]  (.D(n_0_676), .CK(n_0_8), .Q(
      baseReadAdress[11]), .QN());
   DFF_X1 \baseReadAdress_reg[10]  (.D(n_0_675), .CK(n_0_8), .Q(
      baseReadAdress[10]), .QN());
   DFF_X1 \baseReadAdress_reg[9]  (.D(n_0_674), .CK(n_0_8), .Q(baseReadAdress[9]), 
      .QN());
   DFF_X1 \baseReadAdress_reg[8]  (.D(n_0_673), .CK(n_0_8), .Q(baseReadAdress[8]), 
      .QN());
   DFF_X1 \baseReadAdress_reg[7]  (.D(n_0_672), .CK(n_0_8), .Q(baseReadAdress[7]), 
      .QN());
   DFF_X1 \baseReadAdress_reg[6]  (.D(n_0_671), .CK(n_0_8), .Q(baseReadAdress[6]), 
      .QN());
   DFF_X1 \baseReadAdress_reg[5]  (.D(n_0_670), .CK(n_0_8), .Q(baseReadAdress[5]), 
      .QN());
   DFF_X1 \baseReadAdress_reg[4]  (.D(n_0_669), .CK(n_0_8), .Q(baseReadAdress[4]), 
      .QN());
   DFF_X1 \baseReadAdress_reg[3]  (.D(n_0_668), .CK(n_0_8), .Q(baseReadAdress[3]), 
      .QN());
   DFF_X1 \baseReadAdress_reg[2]  (.D(n_0_667), .CK(n_0_8), .Q(baseReadAdress[2]), 
      .QN());
   DFF_X1 \baseReadAdress_reg[1]  (.D(n_0_666), .CK(n_0_8), .Q(baseReadAdress[1]), 
      .QN());
   DFF_X1 \baseReadAdress_reg[0]  (.D(n_0_665), .CK(n_0_8), .Q(baseReadAdress[0]), 
      .QN());
   CLKGATETST_X1 clk_gate_kernelCounter_reg (.CK(clk), .E(n_0_442), .SE(1'b0), 
      .GCK(n_0_9));
   DFF_X1 \kernelCounter_reg[31]  (.D(n_0_439), .CK(n_0_9), .Q(kernelCounter[31]), 
      .QN());
   DFF_X1 \kernelCounter_reg[30]  (.D(n_0_362), .CK(n_0_9), .Q(kernelCounter[30]), 
      .QN());
   DFF_X1 \kernelCounter_reg[29]  (.D(n_0_361), .CK(n_0_9), .Q(kernelCounter[29]), 
      .QN());
   DFF_X1 \kernelCounter_reg[28]  (.D(n_0_360), .CK(n_0_9), .Q(kernelCounter[28]), 
      .QN());
   DFF_X1 \kernelCounter_reg[27]  (.D(n_0_359), .CK(n_0_9), .Q(kernelCounter[27]), 
      .QN());
   DFF_X1 \kernelCounter_reg[26]  (.D(n_0_358), .CK(n_0_9), .Q(kernelCounter[26]), 
      .QN());
   DFF_X1 \kernelCounter_reg[25]  (.D(n_0_357), .CK(n_0_9), .Q(kernelCounter[25]), 
      .QN());
   DFF_X1 \kernelCounter_reg[24]  (.D(n_0_356), .CK(n_0_9), .Q(kernelCounter[24]), 
      .QN());
   DFF_X1 \kernelCounter_reg[23]  (.D(n_0_355), .CK(n_0_9), .Q(kernelCounter[23]), 
      .QN());
   DFF_X1 \kernelCounter_reg[22]  (.D(n_0_354), .CK(n_0_9), .Q(kernelCounter[22]), 
      .QN());
   DFF_X1 \kernelCounter_reg[21]  (.D(n_0_353), .CK(n_0_9), .Q(kernelCounter[21]), 
      .QN());
   DFF_X1 \kernelCounter_reg[20]  (.D(n_0_352), .CK(n_0_9), .Q(kernelCounter[20]), 
      .QN());
   DFF_X1 \kernelCounter_reg[19]  (.D(n_0_351), .CK(n_0_9), .Q(kernelCounter[19]), 
      .QN());
   DFF_X1 \kernelCounter_reg[18]  (.D(n_0_350), .CK(n_0_9), .Q(kernelCounter[18]), 
      .QN());
   DFF_X1 \kernelCounter_reg[17]  (.D(n_0_349), .CK(n_0_9), .Q(kernelCounter[17]), 
      .QN());
   DFF_X1 \kernelCounter_reg[16]  (.D(n_0_348), .CK(n_0_9), .Q(kernelCounter[16]), 
      .QN());
   DFF_X1 \kernelCounter_reg[15]  (.D(n_0_347), .CK(n_0_9), .Q(kernelCounter[15]), 
      .QN());
   DFF_X1 \kernelCounter_reg[14]  (.D(n_0_346), .CK(n_0_9), .Q(kernelCounter[14]), 
      .QN());
   DFF_X1 \kernelCounter_reg[13]  (.D(n_0_345), .CK(n_0_9), .Q(kernelCounter[13]), 
      .QN());
   DFF_X1 \kernelCounter_reg[12]  (.D(n_0_344), .CK(n_0_9), .Q(kernelCounter[12]), 
      .QN());
   DFF_X1 \kernelCounter_reg[11]  (.D(n_0_294), .CK(n_0_9), .Q(kernelCounter[11]), 
      .QN());
   DFF_X1 \kernelCounter_reg[10]  (.D(n_0_293), .CK(n_0_9), .Q(kernelCounter[10]), 
      .QN());
   DFF_X1 \kernelCounter_reg[9]  (.D(n_0_292), .CK(n_0_9), .Q(kernelCounter[9]), 
      .QN());
   DFF_X1 \kernelCounter_reg[8]  (.D(n_0_291), .CK(n_0_9), .Q(kernelCounter[8]), 
      .QN());
   DFF_X1 \kernelCounter_reg[7]  (.D(n_0_290), .CK(n_0_9), .Q(kernelCounter[7]), 
      .QN());
   DFF_X1 \kernelCounter_reg[6]  (.D(n_0_289), .CK(n_0_9), .Q(kernelCounter[6]), 
      .QN());
   DFF_X1 \kernelCounter_reg[5]  (.D(n_0_288), .CK(n_0_9), .Q(kernelCounter[5]), 
      .QN());
   DFF_X1 \kernelCounter_reg[4]  (.D(n_0_287), .CK(n_0_9), .Q(kernelCounter[4]), 
      .QN());
   DFF_X1 \kernelCounter_reg[3]  (.D(n_0_286), .CK(n_0_9), .Q(kernelCounter[3]), 
      .QN());
   DFF_X1 \kernelCounter_reg[2]  (.D(n_0_285), .CK(n_0_9), .Q(kernelCounter[2]), 
      .QN());
   DFF_X1 \kernelCounter_reg[1]  (.D(n_0_284), .CK(n_0_9), .Q(kernelCounter[1]), 
      .QN());
   DFF_X1 \kernelCounter_reg[0]  (.D(n_0_283), .CK(n_0_9), .Q(kernelCounter[0]), 
      .QN());
   DFF_X1 \filterCounter_reg[31]  (.D(n_0_524), .CK(n_0_23), .Q(
      filterCounter[31]), .QN());
   DFF_X1 \filterCounter_reg[30]  (.D(n_0_523), .CK(n_0_23), .Q(
      filterCounter[30]), .QN());
   DFF_X1 \filterCounter_reg[29]  (.D(n_0_522), .CK(n_0_23), .Q(
      filterCounter[29]), .QN());
   DFF_X1 \filterCounter_reg[28]  (.D(n_0_521), .CK(n_0_23), .Q(
      filterCounter[28]), .QN());
   DFF_X1 \filterCounter_reg[27]  (.D(n_0_520), .CK(n_0_23), .Q(
      filterCounter[27]), .QN());
   DFF_X1 \filterCounter_reg[26]  (.D(n_0_519), .CK(n_0_23), .Q(
      filterCounter[26]), .QN());
   DFF_X1 \filterCounter_reg[25]  (.D(n_0_518), .CK(n_0_23), .Q(
      filterCounter[25]), .QN());
   DFF_X1 \filterCounter_reg[24]  (.D(n_0_517), .CK(n_0_23), .Q(
      filterCounter[24]), .QN());
   DFF_X1 \filterCounter_reg[23]  (.D(n_0_516), .CK(n_0_23), .Q(
      filterCounter[23]), .QN());
   DFF_X1 \filterCounter_reg[22]  (.D(n_0_515), .CK(n_0_23), .Q(
      filterCounter[22]), .QN());
   DFF_X1 \filterCounter_reg[21]  (.D(n_0_514), .CK(n_0_23), .Q(
      filterCounter[21]), .QN());
   DFF_X1 \filterCounter_reg[20]  (.D(n_0_513), .CK(n_0_23), .Q(
      filterCounter[20]), .QN());
   DFF_X1 \filterCounter_reg[19]  (.D(n_0_512), .CK(n_0_23), .Q(
      filterCounter[19]), .QN());
   DFF_X1 \filterCounter_reg[18]  (.D(n_0_511), .CK(n_0_23), .Q(
      filterCounter[18]), .QN());
   DFF_X1 \filterCounter_reg[17]  (.D(n_0_509), .CK(n_0_23), .Q(
      filterCounter[17]), .QN());
   DFF_X1 \filterCounter_reg[16]  (.D(n_0_508), .CK(n_0_23), .Q(
      filterCounter[16]), .QN());
   DFF_X1 \filterCounter_reg[15]  (.D(n_0_507), .CK(n_0_23), .Q(
      filterCounter[15]), .QN());
   DFF_X1 \filterCounter_reg[14]  (.D(n_0_506), .CK(n_0_23), .Q(
      filterCounter[14]), .QN());
   DFF_X1 \filterCounter_reg[13]  (.D(n_0_505), .CK(n_0_23), .Q(
      filterCounter[13]), .QN());
   DFF_X1 \filterCounter_reg[12]  (.D(n_0_24), .CK(n_0_23), .Q(filterCounter[12]), 
      .QN());
   DFF_X1 \filterCounter_reg[11]  (.D(n_0_22), .CK(n_0_23), .Q(filterCounter[11]), 
      .QN());
   DFF_X1 \filterCounter_reg[10]  (.D(n_0_21), .CK(n_0_23), .Q(filterCounter[10]), 
      .QN());
   DFF_X1 \filterCounter_reg[9]  (.D(n_0_20), .CK(n_0_23), .Q(filterCounter[9]), 
      .QN());
   DFF_X1 \filterCounter_reg[8]  (.D(n_0_19), .CK(n_0_23), .Q(filterCounter[8]), 
      .QN());
   DFF_X1 \filterCounter_reg[7]  (.D(n_0_18), .CK(n_0_23), .Q(filterCounter[7]), 
      .QN());
   DFF_X1 \filterCounter_reg[6]  (.D(n_0_17), .CK(n_0_23), .Q(filterCounter[6]), 
      .QN());
   DFF_X1 \filterCounter_reg[5]  (.D(n_0_13), .CK(n_0_23), .Q(filterCounter[5]), 
      .QN());
   DFF_X1 \filterCounter_reg[4]  (.D(n_0_12), .CK(n_0_23), .Q(filterCounter[4]), 
      .QN());
   DFF_X1 \filterCounter_reg[3]  (.D(n_0_11), .CK(n_0_23), .Q(filterCounter[3]), 
      .QN());
   DFF_X1 \filterCounter_reg[2]  (.D(n_0_10), .CK(n_0_23), .Q(filterCounter[2]), 
      .QN());
   DFF_X1 \filterCounter_reg[1]  (.D(n_0_4), .CK(n_0_23), .Q(filterCounter[1]), 
      .QN());
   DFF_X1 \filterCounter_reg[0]  (.D(n_0_0), .CK(n_0_23), .Q(filterCounter[0]), 
      .QN());
   CLKGATETST_X1 clk_gate_convWindowX_reg (.CK(clk), .E(n_0_504), .SE(1'b0), 
      .GCK(n_0_14));
   DFF_X1 \convWindowX_reg[31]  (.D(n_0_503), .CK(n_0_14), .Q(convWindowX[31]), 
      .QN());
   DFF_X1 \convWindowX_reg[30]  (.D(n_0_502), .CK(n_0_14), .Q(convWindowX[30]), 
      .QN());
   DFF_X1 \convWindowX_reg[29]  (.D(n_0_501), .CK(n_0_14), .Q(convWindowX[29]), 
      .QN());
   DFF_X1 \convWindowX_reg[28]  (.D(n_0_500), .CK(n_0_14), .Q(convWindowX[28]), 
      .QN());
   DFF_X1 \convWindowX_reg[27]  (.D(n_0_499), .CK(n_0_14), .Q(convWindowX[27]), 
      .QN());
   DFF_X1 \convWindowX_reg[26]  (.D(n_0_498), .CK(n_0_14), .Q(convWindowX[26]), 
      .QN());
   DFF_X1 \convWindowX_reg[25]  (.D(n_0_497), .CK(n_0_14), .Q(convWindowX[25]), 
      .QN());
   DFF_X1 \convWindowX_reg[24]  (.D(n_0_496), .CK(n_0_14), .Q(convWindowX[24]), 
      .QN());
   DFF_X1 \convWindowX_reg[23]  (.D(n_0_495), .CK(n_0_14), .Q(convWindowX[23]), 
      .QN());
   DFF_X1 \convWindowX_reg[22]  (.D(n_0_494), .CK(n_0_14), .Q(convWindowX[22]), 
      .QN());
   DFF_X1 \convWindowX_reg[21]  (.D(n_0_493), .CK(n_0_14), .Q(convWindowX[21]), 
      .QN());
   DFF_X1 \convWindowX_reg[20]  (.D(n_0_492), .CK(n_0_14), .Q(convWindowX[20]), 
      .QN());
   DFF_X1 \convWindowX_reg[19]  (.D(n_0_491), .CK(n_0_14), .Q(convWindowX[19]), 
      .QN());
   DFF_X1 \convWindowX_reg[18]  (.D(n_0_490), .CK(n_0_14), .Q(convWindowX[18]), 
      .QN());
   DFF_X1 \convWindowX_reg[17]  (.D(n_0_489), .CK(n_0_14), .Q(convWindowX[17]), 
      .QN());
   DFF_X1 \convWindowX_reg[16]  (.D(n_0_488), .CK(n_0_14), .Q(convWindowX[16]), 
      .QN());
   DFF_X1 \convWindowX_reg[15]  (.D(n_0_487), .CK(n_0_14), .Q(convWindowX[15]), 
      .QN());
   DFF_X1 \convWindowX_reg[14]  (.D(n_0_457), .CK(n_0_14), .Q(convWindowX[14]), 
      .QN());
   DFF_X1 \convWindowX_reg[13]  (.D(n_0_456), .CK(n_0_14), .Q(convWindowX[13]), 
      .QN());
   DFF_X1 \convWindowX_reg[12]  (.D(n_0_455), .CK(n_0_14), .Q(convWindowX[12]), 
      .QN());
   DFF_X1 \convWindowX_reg[11]  (.D(n_0_454), .CK(n_0_14), .Q(convWindowX[11]), 
      .QN());
   DFF_X1 \convWindowX_reg[10]  (.D(n_0_453), .CK(n_0_14), .Q(convWindowX[10]), 
      .QN());
   DFF_X1 \convWindowX_reg[9]  (.D(n_0_452), .CK(n_0_14), .Q(convWindowX[9]), 
      .QN());
   DFF_X1 \convWindowX_reg[8]  (.D(n_0_451), .CK(n_0_14), .Q(convWindowX[8]), 
      .QN());
   DFF_X1 \convWindowX_reg[7]  (.D(n_0_450), .CK(n_0_14), .Q(convWindowX[7]), 
      .QN());
   DFF_X1 \convWindowX_reg[6]  (.D(n_0_449), .CK(n_0_14), .Q(convWindowX[6]), 
      .QN());
   DFF_X1 \convWindowX_reg[5]  (.D(n_0_448), .CK(n_0_14), .Q(convWindowX[5]), 
      .QN());
   DFF_X1 \convWindowX_reg[4]  (.D(n_0_447), .CK(n_0_14), .Q(convWindowX[4]), 
      .QN());
   DFF_X1 \convWindowX_reg[3]  (.D(n_0_446), .CK(n_0_14), .Q(convWindowX[3]), 
      .QN());
   DFF_X1 \convWindowX_reg[2]  (.D(n_0_445), .CK(n_0_14), .Q(convWindowX[2]), 
      .QN());
   DFF_X1 \convWindowX_reg[1]  (.D(n_0_444), .CK(n_0_14), .Q(convWindowX[1]), 
      .QN());
   DFF_X1 \convWindowX_reg[0]  (.D(n_0_443), .CK(n_0_14), .Q(convWindowX[0]), 
      .QN());
   CLKGATETST_X1 clk_gate_poolingCounter_reg (.CK(clk), .E(n_0_148), .SE(1'b0), 
      .GCK(n_0_15));
   DFF_X1 \poolingCounter_reg[31]  (.D(n_0_147), .CK(n_0_15), .Q(
      poolingCounter[31]), .QN());
   DFF_X1 \poolingCounter_reg[30]  (.D(n_0_146), .CK(n_0_15), .Q(
      poolingCounter[30]), .QN());
   DFF_X1 \poolingCounter_reg[29]  (.D(n_0_145), .CK(n_0_15), .Q(
      poolingCounter[29]), .QN());
   DFF_X1 \poolingCounter_reg[28]  (.D(n_0_144), .CK(n_0_15), .Q(
      poolingCounter[28]), .QN());
   DFF_X1 \poolingCounter_reg[27]  (.D(n_0_143), .CK(n_0_15), .Q(
      poolingCounter[27]), .QN());
   DFF_X1 \poolingCounter_reg[26]  (.D(n_0_142), .CK(n_0_15), .Q(
      poolingCounter[26]), .QN());
   DFF_X1 \poolingCounter_reg[25]  (.D(n_0_141), .CK(n_0_15), .Q(
      poolingCounter[25]), .QN());
   DFF_X1 \poolingCounter_reg[24]  (.D(n_0_140), .CK(n_0_15), .Q(
      poolingCounter[24]), .QN());
   DFF_X1 \poolingCounter_reg[23]  (.D(n_0_139), .CK(n_0_15), .Q(
      poolingCounter[23]), .QN());
   DFF_X1 \poolingCounter_reg[22]  (.D(n_0_138), .CK(n_0_15), .Q(
      poolingCounter[22]), .QN());
   DFF_X1 \poolingCounter_reg[21]  (.D(n_0_137), .CK(n_0_15), .Q(
      poolingCounter[21]), .QN());
   DFF_X1 \poolingCounter_reg[20]  (.D(n_0_129), .CK(n_0_15), .Q(
      poolingCounter[20]), .QN());
   DFF_X1 \poolingCounter_reg[19]  (.D(n_0_128), .CK(n_0_15), .Q(
      poolingCounter[19]), .QN());
   DFF_X1 \poolingCounter_reg[18]  (.D(n_0_127), .CK(n_0_15), .Q(
      poolingCounter[18]), .QN());
   DFF_X1 \poolingCounter_reg[17]  (.D(n_0_126), .CK(n_0_15), .Q(
      poolingCounter[17]), .QN());
   DFF_X1 \poolingCounter_reg[16]  (.D(n_0_125), .CK(n_0_15), .Q(
      poolingCounter[16]), .QN());
   DFF_X1 \poolingCounter_reg[15]  (.D(n_0_124), .CK(n_0_15), .Q(
      poolingCounter[15]), .QN());
   DFF_X1 \poolingCounter_reg[14]  (.D(n_0_123), .CK(n_0_15), .Q(
      poolingCounter[14]), .QN());
   DFF_X1 \poolingCounter_reg[13]  (.D(n_0_122), .CK(n_0_15), .Q(
      poolingCounter[13]), .QN());
   DFF_X1 \poolingCounter_reg[12]  (.D(n_0_121), .CK(n_0_15), .Q(
      poolingCounter[12]), .QN());
   DFF_X1 \poolingCounter_reg[11]  (.D(n_0_120), .CK(n_0_15), .Q(
      poolingCounter[11]), .QN());
   DFF_X1 \poolingCounter_reg[10]  (.D(n_0_110), .CK(n_0_15), .Q(
      poolingCounter[10]), .QN());
   DFF_X1 \poolingCounter_reg[9]  (.D(n_0_77), .CK(n_0_15), .Q(poolingCounter[9]), 
      .QN());
   DFF_X1 \poolingCounter_reg[8]  (.D(n_0_76), .CK(n_0_15), .Q(poolingCounter[8]), 
      .QN());
   DFF_X1 \poolingCounter_reg[7]  (.D(n_0_75), .CK(n_0_15), .Q(poolingCounter[7]), 
      .QN());
   DFF_X1 \poolingCounter_reg[6]  (.D(n_0_74), .CK(n_0_15), .Q(poolingCounter[6]), 
      .QN());
   DFF_X1 \poolingCounter_reg[5]  (.D(n_0_73), .CK(n_0_15), .Q(poolingCounter[5]), 
      .QN());
   DFF_X1 \poolingCounter_reg[4]  (.D(n_0_72), .CK(n_0_15), .Q(poolingCounter[4]), 
      .QN());
   DFF_X1 \poolingCounter_reg[3]  (.D(n_0_56), .CK(n_0_15), .Q(poolingCounter[3]), 
      .QN());
   DFF_X1 \poolingCounter_reg[2]  (.D(n_0_37), .CK(n_0_15), .Q(poolingCounter[2]), 
      .QN());
   DFF_X1 \poolingCounter_reg[1]  (.D(n_0_35), .CK(n_0_15), .Q(poolingCounter[1]), 
      .QN());
   DFF_X1 \poolingCounter_reg[0]  (.D(n_0_33), .CK(n_0_15), .Q(poolingCounter[0]), 
      .QN());
   CLKGATETST_X1 clk_gate_poolingWindowX_reg (.CK(clk), .E(n_0_199), .SE(1'b0), 
      .GCK(n_0_16));
   DFF_X1 \poolingWindowX_reg[31]  (.D(n_0_198), .CK(n_0_16), .Q(
      poolingWindowX[31]), .QN());
   DFF_X1 \poolingWindowX_reg[30]  (.D(n_0_197), .CK(n_0_16), .Q(
      poolingWindowX[30]), .QN());
   DFF_X1 \poolingWindowX_reg[29]  (.D(n_0_196), .CK(n_0_16), .Q(
      poolingWindowX[29]), .QN());
   DFF_X1 \poolingWindowX_reg[28]  (.D(n_0_195), .CK(n_0_16), .Q(
      poolingWindowX[28]), .QN());
   DFF_X1 \poolingWindowX_reg[27]  (.D(n_0_194), .CK(n_0_16), .Q(
      poolingWindowX[27]), .QN());
   DFF_X1 \poolingWindowX_reg[26]  (.D(n_0_193), .CK(n_0_16), .Q(
      poolingWindowX[26]), .QN());
   DFF_X1 \poolingWindowX_reg[25]  (.D(n_0_192), .CK(n_0_16), .Q(
      poolingWindowX[25]), .QN());
   DFF_X1 \poolingWindowX_reg[24]  (.D(n_0_191), .CK(n_0_16), .Q(
      poolingWindowX[24]), .QN());
   DFF_X1 \poolingWindowX_reg[23]  (.D(n_0_190), .CK(n_0_16), .Q(
      poolingWindowX[23]), .QN());
   DFF_X1 \poolingWindowX_reg[22]  (.D(n_0_189), .CK(n_0_16), .Q(
      poolingWindowX[22]), .QN());
   DFF_X1 \poolingWindowX_reg[21]  (.D(n_0_188), .CK(n_0_16), .Q(
      poolingWindowX[21]), .QN());
   DFF_X1 \poolingWindowX_reg[20]  (.D(n_0_187), .CK(n_0_16), .Q(
      poolingWindowX[20]), .QN());
   DFF_X1 \poolingWindowX_reg[19]  (.D(n_0_186), .CK(n_0_16), .Q(
      poolingWindowX[19]), .QN());
   DFF_X1 \poolingWindowX_reg[18]  (.D(n_0_185), .CK(n_0_16), .Q(
      poolingWindowX[18]), .QN());
   DFF_X1 \poolingWindowX_reg[17]  (.D(n_0_184), .CK(n_0_16), .Q(
      poolingWindowX[17]), .QN());
   DFF_X1 \poolingWindowX_reg[16]  (.D(n_0_164), .CK(n_0_16), .Q(
      poolingWindowX[16]), .QN());
   DFF_X1 \poolingWindowX_reg[15]  (.D(n_0_163), .CK(n_0_16), .Q(
      poolingWindowX[15]), .QN());
   DFF_X1 \poolingWindowX_reg[14]  (.D(n_0_162), .CK(n_0_16), .Q(
      poolingWindowX[14]), .QN());
   DFF_X1 \poolingWindowX_reg[13]  (.D(n_0_161), .CK(n_0_16), .Q(
      poolingWindowX[13]), .QN());
   DFF_X1 \poolingWindowX_reg[12]  (.D(n_0_160), .CK(n_0_16), .Q(
      poolingWindowX[12]), .QN());
   DFF_X1 \poolingWindowX_reg[11]  (.D(n_0_159), .CK(n_0_16), .Q(
      poolingWindowX[11]), .QN());
   DFF_X1 \poolingWindowX_reg[10]  (.D(n_0_158), .CK(n_0_16), .Q(
      poolingWindowX[10]), .QN());
   DFF_X1 \poolingWindowX_reg[9]  (.D(n_0_157), .CK(n_0_16), .Q(
      poolingWindowX[9]), .QN());
   DFF_X1 \poolingWindowX_reg[8]  (.D(n_0_156), .CK(n_0_16), .Q(
      poolingWindowX[8]), .QN());
   DFF_X1 \poolingWindowX_reg[7]  (.D(n_0_155), .CK(n_0_16), .Q(
      poolingWindowX[7]), .QN());
   DFF_X1 \poolingWindowX_reg[6]  (.D(n_0_154), .CK(n_0_16), .Q(
      poolingWindowX[6]), .QN());
   DFF_X1 \poolingWindowX_reg[5]  (.D(n_0_153), .CK(n_0_16), .Q(
      poolingWindowX[5]), .QN());
   DFF_X1 \poolingWindowX_reg[4]  (.D(n_0_152), .CK(n_0_16), .Q(
      poolingWindowX[4]), .QN());
   DFF_X1 \poolingWindowX_reg[3]  (.D(n_0_151), .CK(n_0_16), .Q(
      poolingWindowX[3]), .QN());
   DFF_X1 \poolingWindowX_reg[2]  (.D(n_0_150), .CK(n_0_16), .Q(
      poolingWindowX[2]), .QN());
   DFF_X1 \poolingWindowX_reg[1]  (.D(n_0_149), .CK(n_0_16), .Q(
      poolingWindowX[1]), .QN());
   CLKGATETST_X1 clk_gate_poolingWindowY_reg (.CK(clk), .E(n_0_275), .SE(1'b0), 
      .GCK(n_0_510));
   DFF_X1 \poolingWindowY_reg[31]  (.D(n_0_274), .CK(n_0_510), .Q(
      poolingWindowY[31]), .QN());
   DFF_X1 \poolingWindowY_reg[30]  (.D(n_0_273), .CK(n_0_510), .Q(
      poolingWindowY[30]), .QN());
   DFF_X1 \poolingWindowY_reg[29]  (.D(n_0_272), .CK(n_0_510), .Q(
      poolingWindowY[29]), .QN());
   DFF_X1 \poolingWindowY_reg[28]  (.D(n_0_271), .CK(n_0_510), .Q(
      poolingWindowY[28]), .QN());
   DFF_X1 \poolingWindowY_reg[27]  (.D(n_0_270), .CK(n_0_510), .Q(
      poolingWindowY[27]), .QN());
   DFF_X1 \poolingWindowY_reg[26]  (.D(n_0_269), .CK(n_0_510), .Q(
      poolingWindowY[26]), .QN());
   DFF_X1 \poolingWindowY_reg[25]  (.D(n_0_268), .CK(n_0_510), .Q(
      poolingWindowY[25]), .QN());
   DFF_X1 \poolingWindowY_reg[24]  (.D(n_0_267), .CK(n_0_510), .Q(
      poolingWindowY[24]), .QN());
   DFF_X1 \poolingWindowY_reg[23]  (.D(n_0_266), .CK(n_0_510), .Q(
      poolingWindowY[23]), .QN());
   DFF_X1 \poolingWindowY_reg[22]  (.D(n_0_265), .CK(n_0_510), .Q(
      poolingWindowY[22]), .QN());
   DFF_X1 \poolingWindowY_reg[21]  (.D(n_0_264), .CK(n_0_510), .Q(
      poolingWindowY[21]), .QN());
   DFF_X1 \poolingWindowY_reg[20]  (.D(n_0_263), .CK(n_0_510), .Q(
      poolingWindowY[20]), .QN());
   DFF_X1 \poolingWindowY_reg[19]  (.D(n_0_262), .CK(n_0_510), .Q(
      poolingWindowY[19]), .QN());
   DFF_X1 \poolingWindowY_reg[18]  (.D(n_0_234), .CK(n_0_510), .Q(
      poolingWindowY[18]), .QN());
   DFF_X1 \poolingWindowY_reg[17]  (.D(n_0_229), .CK(n_0_510), .Q(
      poolingWindowY[17]), .QN());
   DFF_X1 \poolingWindowY_reg[16]  (.D(n_0_228), .CK(n_0_510), .Q(
      poolingWindowY[16]), .QN());
   DFF_X1 \poolingWindowY_reg[15]  (.D(n_0_227), .CK(n_0_510), .Q(
      poolingWindowY[15]), .QN());
   DFF_X1 \poolingWindowY_reg[14]  (.D(n_0_226), .CK(n_0_510), .Q(
      poolingWindowY[14]), .QN());
   DFF_X1 \poolingWindowY_reg[13]  (.D(n_0_225), .CK(n_0_510), .Q(
      poolingWindowY[13]), .QN());
   DFF_X1 \poolingWindowY_reg[12]  (.D(n_0_224), .CK(n_0_510), .Q(
      poolingWindowY[12]), .QN());
   DFF_X1 \poolingWindowY_reg[11]  (.D(n_0_223), .CK(n_0_510), .Q(
      poolingWindowY[11]), .QN());
   DFF_X1 \poolingWindowY_reg[10]  (.D(n_0_222), .CK(n_0_510), .Q(
      poolingWindowY[10]), .QN());
   DFF_X1 \poolingWindowY_reg[9]  (.D(n_0_221), .CK(n_0_510), .Q(
      poolingWindowY[9]), .QN());
   DFF_X1 \poolingWindowY_reg[8]  (.D(n_0_220), .CK(n_0_510), .Q(
      poolingWindowY[8]), .QN());
   DFF_X1 \poolingWindowY_reg[7]  (.D(n_0_219), .CK(n_0_510), .Q(
      poolingWindowY[7]), .QN());
   DFF_X1 \poolingWindowY_reg[6]  (.D(n_0_218), .CK(n_0_510), .Q(
      poolingWindowY[6]), .QN());
   DFF_X1 \poolingWindowY_reg[5]  (.D(n_0_217), .CK(n_0_510), .Q(
      poolingWindowY[5]), .QN());
   DFF_X1 \poolingWindowY_reg[4]  (.D(n_0_216), .CK(n_0_510), .Q(
      poolingWindowY[4]), .QN());
   DFF_X1 \poolingWindowY_reg[3]  (.D(n_0_215), .CK(n_0_510), .Q(
      poolingWindowY[3]), .QN());
   DFF_X1 \poolingWindowY_reg[2]  (.D(n_0_214), .CK(n_0_510), .Q(
      poolingWindowY[2]), .QN());
   DFF_X1 \poolingWindowY_reg[1]  (.D(n_0_213), .CK(n_0_510), .Q(
      poolingWindowY[1]), .QN());
   CLKGATETST_X1 clk_gate_index_filter_reg (.CK(clk), .E(n_0_36), .SE(1'b0), 
      .GCK(n_0_23));
   HA_X1 i_0_0_678 (.A(layerCounter[2]), .B(n_0_0_65), .CO(n_0_0_1), .S());
   HA_X1 i_0_0_723 (.A(n_0_683), .B(n_0_682), .CO(n_0_0_0), .S(n_0_0_31));
   HA_X1 i_0_0_724 (.A(n_0_684), .B(n_0_0_0), .CO(n_0_0_2), .S(n_0_0_32));
   HA_X1 i_0_0_725 (.A(n_0_685), .B(n_0_0_2), .CO(n_0_0_3), .S(n_0_0_33));
   HA_X1 i_0_0_726 (.A(n_0_686), .B(n_0_0_3), .CO(n_0_0_4), .S(n_0_0_34));
   HA_X1 i_0_0_727 (.A(n_0_687), .B(n_0_0_4), .CO(n_0_0_5), .S(n_0_0_35));
   HA_X1 i_0_0_728 (.A(n_0_688), .B(n_0_0_5), .CO(n_0_0_6), .S(n_0_0_36));
   HA_X1 i_0_0_729 (.A(n_0_689), .B(n_0_0_6), .CO(n_0_0_7), .S(n_0_0_37));
   HA_X1 i_0_0_730 (.A(n_0_690), .B(n_0_0_7), .CO(n_0_0_8), .S(n_0_0_38));
   HA_X1 i_0_0_731 (.A(n_0_691), .B(n_0_0_8), .CO(n_0_0_9), .S(n_0_0_39));
   HA_X1 i_0_0_732 (.A(n_0_692), .B(n_0_0_9), .CO(n_0_0_10), .S(n_0_0_40));
   HA_X1 i_0_0_733 (.A(n_0_693), .B(n_0_0_10), .CO(n_0_0_11), .S(n_0_0_41));
   HA_X1 i_0_0_734 (.A(n_0_694), .B(n_0_0_11), .CO(n_0_0_12), .S(n_0_0_42));
   HA_X1 i_0_0_735 (.A(n_0_695), .B(n_0_0_12), .CO(n_0_0_13), .S(n_0_0_43));
   FA_X1 i_0_0_798 (.A(1'b0), .B(n_0_548), .CI(n_0_571), .CO(n_0_0_59), .S(
      n_0_639));
   FA_X1 i_0_0_799 (.A(n_0_0_62), .B(n_0_646), .CI(n_0_0_59), .CO(n_0_0_60), 
      .S(n_0_640));
   FA_X1 i_0_0_800 (.A(1'b0), .B(n_0_581), .CI(n_0_0_60), .CO(n_0_642), .S(
      n_0_641));
   FA_X1 i_0_0_845 (.A(n_0_540), .B(n_0_0_61), .CI(n_0_539), .CO(n_0_0_14), 
      .S(n_0_0_44));
   FA_X1 i_0_0_846 (.A(n_0_541), .B(n_0_0_28), .CI(n_0_0_14), .CO(n_0_0_15), 
      .S(n_0_0_45));
   FA_X1 i_0_0_847 (.A(n_0_542), .B(n_0_0_29), .CI(n_0_0_15), .CO(n_0_0_16), 
      .S(n_0_0_46));
   FA_X1 i_0_0_848 (.A(n_0_543), .B(n_0_0_30), .CI(n_0_0_16), .CO(n_0_0_17), 
      .S(n_0_0_47));
   FA_X1 i_0_0_849 (.A(n_0_544), .B(n_0_0_55), .CI(n_0_0_17), .CO(n_0_0_18), 
      .S(n_0_0_48));
   FA_X1 i_0_0_850 (.A(n_0_545), .B(n_0_572), .CI(n_0_0_18), .CO(n_0_0_19), 
      .S(n_0_0_49));
   FA_X1 i_0_0_851 (.A(n_0_546), .B(n_0_0_56), .CI(n_0_0_19), .CO(n_0_0_20), 
      .S(n_0_0_50));
   FA_X1 i_0_0_852 (.A(n_0_0_57), .B(n_0_547), .CI(n_0_0_20), .CO(n_0_0_21), 
      .S(n_0_0_51));
   FA_X1 i_0_0_853 (.A(n_0_0_27), .B(n_0_0_58), .CI(n_0_0_21), .CO(n_0_0_22), 
      .S(n_0_0_52));
   FA_X1 i_0_0_854 (.A(n_0_571), .B(n_0_0_58), .CI(n_0_0_22), .CO(n_0_0_23), 
      .S(n_0_0_53));
   FA_X1 i_0_0_855 (.A(n_0_0_61), .B(n_0_0_58), .CI(n_0_0_23), .CO(n_0_0_24), 
      .S(n_0_0_54));
   HA_X1 i_0_0_888 (.A(layerCounter[1]), .B(layerCounter[0]), .CO(n_0_0_25), 
      .S(n_0_0_63));
   HA_X1 i_0_0_889 (.A(layerCounter[2]), .B(n_0_0_25), .CO(n_0_0_26), .S(
      n_0_0_64));
   OAI22_X1 i_0_0_14 (.A1(n_0_0_81), .A2(n_0_0_75), .B1(n_0_0_80), .B2(n_0_0_431), 
      .ZN(n_0_550));
   NOR2_X1 i_0_0_15 (.A1(n_0_0_431), .A2(n_0_0_71), .ZN(n_0_0_75));
   NOR2_X1 i_0_0_16 (.A1(layerCounter[0]), .A2(reset), .ZN(n_0_26));
   AND2_X1 i_0_0_17 (.A1(n_0_0_73), .A2(n_0_0_63), .ZN(n_0_27));
   AND2_X1 i_0_0_18 (.A1(n_0_0_73), .A2(n_0_0_64), .ZN(n_0_28));
   NOR2_X1 i_0_0_19 (.A1(reset), .A2(n_0_0_77), .ZN(n_0_29));
   XNOR2_X1 i_0_0_20 (.A(layerCounter[31]), .B(n_0_0_26), .ZN(n_0_0_77));
   NOR2_X1 i_0_0_21 (.A1(n_0_0_209), .A2(poolingCounter[0]), .ZN(n_0_33));
   AND2_X1 i_0_0_22 (.A1(n_0_440), .A2(n_0_563), .ZN(n_0_35));
   AND2_X1 i_0_0_23 (.A1(n_0_441), .A2(n_0_563), .ZN(n_0_37));
   AND2_X1 i_0_0_24 (.A1(n_0_458), .A2(n_0_563), .ZN(n_0_56));
   AND2_X1 i_0_0_25 (.A1(n_0_459), .A2(n_0_563), .ZN(n_0_72));
   AND2_X1 i_0_0_26 (.A1(n_0_460), .A2(n_0_563), .ZN(n_0_73));
   AND2_X1 i_0_0_27 (.A1(n_0_461), .A2(n_0_563), .ZN(n_0_74));
   AND2_X1 i_0_0_28 (.A1(n_0_462), .A2(n_0_563), .ZN(n_0_75));
   AND2_X1 i_0_0_29 (.A1(n_0_463), .A2(n_0_563), .ZN(n_0_76));
   AND2_X1 i_0_0_30 (.A1(n_0_464), .A2(n_0_563), .ZN(n_0_77));
   AND2_X1 i_0_0_31 (.A1(n_0_465), .A2(n_0_563), .ZN(n_0_110));
   AND2_X1 i_0_0_32 (.A1(n_0_466), .A2(n_0_563), .ZN(n_0_120));
   AND2_X1 i_0_0_33 (.A1(n_0_467), .A2(n_0_563), .ZN(n_0_121));
   AND2_X1 i_0_0_34 (.A1(n_0_468), .A2(n_0_563), .ZN(n_0_122));
   AND2_X1 i_0_0_35 (.A1(n_0_469), .A2(n_0_563), .ZN(n_0_123));
   AND2_X1 i_0_0_36 (.A1(n_0_470), .A2(n_0_563), .ZN(n_0_124));
   AND2_X1 i_0_0_37 (.A1(n_0_471), .A2(n_0_563), .ZN(n_0_125));
   AND2_X1 i_0_0_38 (.A1(n_0_472), .A2(n_0_563), .ZN(n_0_126));
   AND2_X1 i_0_0_39 (.A1(n_0_473), .A2(n_0_563), .ZN(n_0_127));
   AND2_X1 i_0_0_40 (.A1(n_0_474), .A2(n_0_563), .ZN(n_0_128));
   AND2_X1 i_0_0_41 (.A1(n_0_475), .A2(n_0_563), .ZN(n_0_129));
   AND2_X1 i_0_0_42 (.A1(n_0_476), .A2(n_0_563), .ZN(n_0_137));
   AND2_X1 i_0_0_43 (.A1(n_0_477), .A2(n_0_563), .ZN(n_0_138));
   AND2_X1 i_0_0_44 (.A1(n_0_478), .A2(n_0_563), .ZN(n_0_139));
   AND2_X1 i_0_0_45 (.A1(n_0_479), .A2(n_0_563), .ZN(n_0_140));
   AND2_X1 i_0_0_46 (.A1(n_0_480), .A2(n_0_563), .ZN(n_0_141));
   AND2_X1 i_0_0_47 (.A1(n_0_481), .A2(n_0_563), .ZN(n_0_142));
   AND2_X1 i_0_0_48 (.A1(n_0_482), .A2(n_0_563), .ZN(n_0_143));
   AND2_X1 i_0_0_49 (.A1(n_0_483), .A2(n_0_563), .ZN(n_0_144));
   AND2_X1 i_0_0_50 (.A1(n_0_484), .A2(n_0_563), .ZN(n_0_145));
   AND2_X1 i_0_0_51 (.A1(n_0_485), .A2(n_0_563), .ZN(n_0_146));
   AND2_X1 i_0_0_52 (.A1(n_0_486), .A2(n_0_563), .ZN(n_0_147));
   NOR2_X1 i_0_0_53 (.A1(n_0_0_210), .A2(n_0_0_78), .ZN(n_0_148));
   AND2_X1 i_0_0_54 (.A1(n_0_408), .A2(n_0_0_78), .ZN(n_0_149));
   AND2_X1 i_0_0_55 (.A1(n_0_409), .A2(n_0_0_78), .ZN(n_0_150));
   AND2_X1 i_0_0_56 (.A1(n_0_410), .A2(n_0_0_78), .ZN(n_0_151));
   AND2_X1 i_0_0_57 (.A1(n_0_411), .A2(n_0_0_78), .ZN(n_0_152));
   AND2_X1 i_0_0_58 (.A1(n_0_412), .A2(n_0_0_78), .ZN(n_0_153));
   AND2_X1 i_0_0_59 (.A1(n_0_413), .A2(n_0_0_78), .ZN(n_0_154));
   AND2_X1 i_0_0_60 (.A1(n_0_414), .A2(n_0_0_78), .ZN(n_0_155));
   AND2_X1 i_0_0_61 (.A1(n_0_415), .A2(n_0_0_78), .ZN(n_0_156));
   AND2_X1 i_0_0_62 (.A1(n_0_416), .A2(n_0_0_78), .ZN(n_0_157));
   AND2_X1 i_0_0_63 (.A1(n_0_417), .A2(n_0_0_78), .ZN(n_0_158));
   AND2_X1 i_0_0_64 (.A1(n_0_418), .A2(n_0_0_78), .ZN(n_0_159));
   AND2_X1 i_0_0_65 (.A1(n_0_419), .A2(n_0_0_78), .ZN(n_0_160));
   AND2_X1 i_0_0_66 (.A1(n_0_420), .A2(n_0_0_78), .ZN(n_0_161));
   AND2_X1 i_0_0_67 (.A1(n_0_421), .A2(n_0_0_78), .ZN(n_0_162));
   AND2_X1 i_0_0_68 (.A1(n_0_422), .A2(n_0_0_78), .ZN(n_0_163));
   AND2_X1 i_0_0_69 (.A1(n_0_423), .A2(n_0_0_78), .ZN(n_0_164));
   AND2_X1 i_0_0_70 (.A1(n_0_424), .A2(n_0_0_78), .ZN(n_0_184));
   AND2_X1 i_0_0_71 (.A1(n_0_425), .A2(n_0_0_78), .ZN(n_0_185));
   AND2_X1 i_0_0_72 (.A1(n_0_426), .A2(n_0_0_78), .ZN(n_0_186));
   AND2_X1 i_0_0_73 (.A1(n_0_427), .A2(n_0_0_78), .ZN(n_0_187));
   AND2_X1 i_0_0_74 (.A1(n_0_428), .A2(n_0_0_78), .ZN(n_0_188));
   AND2_X1 i_0_0_75 (.A1(n_0_429), .A2(n_0_0_78), .ZN(n_0_189));
   AND2_X1 i_0_0_76 (.A1(n_0_430), .A2(n_0_0_78), .ZN(n_0_190));
   AND2_X1 i_0_0_77 (.A1(n_0_431), .A2(n_0_0_78), .ZN(n_0_191));
   AND2_X1 i_0_0_78 (.A1(n_0_432), .A2(n_0_0_78), .ZN(n_0_192));
   AND2_X1 i_0_0_79 (.A1(n_0_433), .A2(n_0_0_78), .ZN(n_0_193));
   AND2_X1 i_0_0_80 (.A1(n_0_434), .A2(n_0_0_78), .ZN(n_0_194));
   AND2_X1 i_0_0_81 (.A1(n_0_435), .A2(n_0_0_78), .ZN(n_0_195));
   AND2_X1 i_0_0_82 (.A1(n_0_436), .A2(n_0_0_78), .ZN(n_0_196));
   AND2_X1 i_0_0_83 (.A1(n_0_437), .A2(n_0_0_78), .ZN(n_0_197));
   AND2_X1 i_0_0_84 (.A1(n_0_438), .A2(n_0_0_78), .ZN(n_0_198));
   NOR2_X1 i_0_0_85 (.A1(n_0_0_209), .A2(n_0_0_328), .ZN(n_0_0_78));
   AOI21_X1 i_0_0_86 (.A(n_0_0_79), .B1(n_0_0_304), .B2(n_0_0_73), .ZN(n_0_199));
   AND2_X1 i_0_0_87 (.A1(n_0_377), .A2(n_0_0_79), .ZN(n_0_213));
   AND2_X1 i_0_0_88 (.A1(n_0_378), .A2(n_0_0_79), .ZN(n_0_214));
   AND2_X1 i_0_0_89 (.A1(n_0_379), .A2(n_0_0_79), .ZN(n_0_215));
   AND2_X1 i_0_0_90 (.A1(n_0_380), .A2(n_0_0_79), .ZN(n_0_216));
   AND2_X1 i_0_0_91 (.A1(n_0_381), .A2(n_0_0_79), .ZN(n_0_217));
   AND2_X1 i_0_0_92 (.A1(n_0_382), .A2(n_0_0_79), .ZN(n_0_218));
   AND2_X1 i_0_0_93 (.A1(n_0_383), .A2(n_0_0_79), .ZN(n_0_219));
   AND2_X1 i_0_0_94 (.A1(n_0_384), .A2(n_0_0_79), .ZN(n_0_220));
   AND2_X1 i_0_0_95 (.A1(n_0_385), .A2(n_0_0_79), .ZN(n_0_221));
   AND2_X1 i_0_0_96 (.A1(n_0_386), .A2(n_0_0_79), .ZN(n_0_222));
   AND2_X1 i_0_0_97 (.A1(n_0_387), .A2(n_0_0_79), .ZN(n_0_223));
   AND2_X1 i_0_0_98 (.A1(n_0_388), .A2(n_0_0_79), .ZN(n_0_224));
   AND2_X1 i_0_0_99 (.A1(n_0_389), .A2(n_0_0_79), .ZN(n_0_225));
   AND2_X1 i_0_0_100 (.A1(n_0_390), .A2(n_0_0_79), .ZN(n_0_226));
   AND2_X1 i_0_0_101 (.A1(n_0_391), .A2(n_0_0_79), .ZN(n_0_227));
   AND2_X1 i_0_0_102 (.A1(n_0_392), .A2(n_0_0_79), .ZN(n_0_228));
   AND2_X1 i_0_0_103 (.A1(n_0_393), .A2(n_0_0_79), .ZN(n_0_229));
   AND2_X1 i_0_0_104 (.A1(n_0_394), .A2(n_0_0_79), .ZN(n_0_234));
   AND2_X1 i_0_0_105 (.A1(n_0_395), .A2(n_0_0_79), .ZN(n_0_262));
   AND2_X1 i_0_0_106 (.A1(n_0_396), .A2(n_0_0_79), .ZN(n_0_263));
   AND2_X1 i_0_0_107 (.A1(n_0_397), .A2(n_0_0_79), .ZN(n_0_264));
   AND2_X1 i_0_0_108 (.A1(n_0_398), .A2(n_0_0_79), .ZN(n_0_265));
   AND2_X1 i_0_0_109 (.A1(n_0_399), .A2(n_0_0_79), .ZN(n_0_266));
   AND2_X1 i_0_0_110 (.A1(n_0_400), .A2(n_0_0_79), .ZN(n_0_267));
   AND2_X1 i_0_0_111 (.A1(n_0_401), .A2(n_0_0_79), .ZN(n_0_268));
   AND2_X1 i_0_0_112 (.A1(n_0_402), .A2(n_0_0_79), .ZN(n_0_269));
   AND2_X1 i_0_0_113 (.A1(n_0_403), .A2(n_0_0_79), .ZN(n_0_270));
   AND2_X1 i_0_0_114 (.A1(n_0_404), .A2(n_0_0_79), .ZN(n_0_271));
   AND2_X1 i_0_0_115 (.A1(n_0_405), .A2(n_0_0_79), .ZN(n_0_272));
   AND2_X1 i_0_0_116 (.A1(n_0_406), .A2(n_0_0_79), .ZN(n_0_273));
   AND2_X1 i_0_0_117 (.A1(n_0_407), .A2(n_0_0_79), .ZN(n_0_274));
   NOR3_X1 i_0_0_118 (.A1(reset), .A2(n_0_0_328), .A3(n_0_0_283), .ZN(n_0_0_79));
   OAI21_X1 i_0_0_119 (.A(n_0_0_73), .B1(n_0_0_303), .B2(n_0_0_281), .ZN(n_0_275));
   NOR2_X1 i_0_0_120 (.A1(n_0_0_278), .A2(n_0_0_84), .ZN(n_0_551));
   INV_X1 i_0_0_121 (.A(n_0_0_80), .ZN(n_0_552));
   NAND3_X1 i_0_0_122 (.A1(n_0_0_73), .A2(n_0_0_71), .A3(poolingState[0]), 
      .ZN(n_0_0_80));
   OAI21_X1 i_0_0_123 (.A(n_0_0_212), .B1(n_0_0_305), .B2(n_0_0_306), .ZN(
      n_0_279));
   OAI22_X1 i_0_0_124 (.A1(n_0_0_428), .A2(n_0_0_84), .B1(n_0_0_81), .B2(
      n_0_0_110), .ZN(n_0_554));
   NAND2_X1 i_0_0_125 (.A1(n_0_0_74), .A2(n_0_0_73), .ZN(n_0_0_81));
   NOR2_X1 i_0_0_126 (.A1(n_0_0_110), .A2(n_0_0_84), .ZN(n_0_555));
   INV_X1 i_0_0_127 (.A(n_0_0_82), .ZN(n_0_556));
   AOI21_X1 i_0_0_128 (.A(reset), .B1(n_0_0_211), .B2(n_0_0_425), .ZN(n_0_0_82));
   AND2_X1 i_0_0_129 (.A1(n_0_326), .A2(n_0_0_215), .ZN(n_0_283));
   AND2_X1 i_0_0_130 (.A1(n_0_327), .A2(n_0_0_215), .ZN(n_0_284));
   AND2_X1 i_0_0_131 (.A1(n_0_328), .A2(n_0_0_215), .ZN(n_0_285));
   AND2_X1 i_0_0_132 (.A1(n_0_329), .A2(n_0_0_215), .ZN(n_0_286));
   AND2_X1 i_0_0_133 (.A1(n_0_330), .A2(n_0_0_215), .ZN(n_0_287));
   AND2_X1 i_0_0_134 (.A1(n_0_331), .A2(n_0_0_215), .ZN(n_0_288));
   AND2_X1 i_0_0_135 (.A1(n_0_332), .A2(n_0_0_215), .ZN(n_0_289));
   AND2_X1 i_0_0_136 (.A1(n_0_333), .A2(n_0_0_215), .ZN(n_0_290));
   AND2_X1 i_0_0_137 (.A1(n_0_334), .A2(n_0_0_215), .ZN(n_0_291));
   AND2_X1 i_0_0_138 (.A1(n_0_335), .A2(n_0_0_215), .ZN(n_0_292));
   AND2_X1 i_0_0_139 (.A1(n_0_336), .A2(n_0_0_215), .ZN(n_0_293));
   AND2_X1 i_0_0_140 (.A1(n_0_337), .A2(n_0_0_215), .ZN(n_0_294));
   AND2_X1 i_0_0_141 (.A1(n_0_338), .A2(n_0_0_215), .ZN(n_0_344));
   AND2_X1 i_0_0_142 (.A1(n_0_339), .A2(n_0_0_215), .ZN(n_0_345));
   AND2_X1 i_0_0_143 (.A1(n_0_340), .A2(n_0_0_215), .ZN(n_0_346));
   AND2_X1 i_0_0_144 (.A1(n_0_341), .A2(n_0_0_215), .ZN(n_0_347));
   AND2_X1 i_0_0_145 (.A1(n_0_342), .A2(n_0_0_215), .ZN(n_0_348));
   AND2_X1 i_0_0_146 (.A1(n_0_343), .A2(n_0_0_215), .ZN(n_0_349));
   AND2_X1 i_0_0_147 (.A1(n_0_363), .A2(n_0_0_215), .ZN(n_0_350));
   AND2_X1 i_0_0_148 (.A1(n_0_364), .A2(n_0_0_215), .ZN(n_0_351));
   AND2_X1 i_0_0_149 (.A1(n_0_365), .A2(n_0_0_215), .ZN(n_0_352));
   AND2_X1 i_0_0_150 (.A1(n_0_366), .A2(n_0_0_215), .ZN(n_0_353));
   AND2_X1 i_0_0_151 (.A1(n_0_367), .A2(n_0_0_215), .ZN(n_0_354));
   AND2_X1 i_0_0_152 (.A1(n_0_368), .A2(n_0_0_215), .ZN(n_0_355));
   AND2_X1 i_0_0_153 (.A1(n_0_369), .A2(n_0_0_215), .ZN(n_0_356));
   AND2_X1 i_0_0_154 (.A1(n_0_370), .A2(n_0_0_215), .ZN(n_0_357));
   AND2_X1 i_0_0_155 (.A1(n_0_371), .A2(n_0_0_215), .ZN(n_0_358));
   AND2_X1 i_0_0_156 (.A1(n_0_372), .A2(n_0_0_215), .ZN(n_0_359));
   AND2_X1 i_0_0_157 (.A1(n_0_373), .A2(n_0_0_215), .ZN(n_0_360));
   AND2_X1 i_0_0_158 (.A1(n_0_374), .A2(n_0_0_215), .ZN(n_0_361));
   AND2_X1 i_0_0_159 (.A1(n_0_375), .A2(n_0_0_215), .ZN(n_0_362));
   AND2_X1 i_0_0_160 (.A1(n_0_376), .A2(n_0_0_215), .ZN(n_0_439));
   NOR2_X1 i_0_0_161 (.A1(n_0_0_213), .A2(n_0_561), .ZN(n_0_442));
   NOR3_X1 i_0_0_162 (.A1(convWindowX[0]), .A2(n_0_0_389), .A3(n_0_0_214), 
      .ZN(n_0_443));
   AND2_X1 i_0_0_163 (.A1(n_0_295), .A2(n_0_561), .ZN(n_0_444));
   AND2_X1 i_0_0_164 (.A1(n_0_296), .A2(n_0_561), .ZN(n_0_445));
   AND2_X1 i_0_0_165 (.A1(n_0_297), .A2(n_0_561), .ZN(n_0_446));
   AND2_X1 i_0_0_166 (.A1(n_0_298), .A2(n_0_561), .ZN(n_0_447));
   AND2_X1 i_0_0_167 (.A1(n_0_299), .A2(n_0_561), .ZN(n_0_448));
   AND2_X1 i_0_0_168 (.A1(n_0_300), .A2(n_0_561), .ZN(n_0_449));
   AND2_X1 i_0_0_169 (.A1(n_0_301), .A2(n_0_561), .ZN(n_0_450));
   AND2_X1 i_0_0_170 (.A1(n_0_302), .A2(n_0_561), .ZN(n_0_451));
   AND2_X1 i_0_0_171 (.A1(n_0_303), .A2(n_0_561), .ZN(n_0_452));
   AND2_X1 i_0_0_172 (.A1(n_0_304), .A2(n_0_561), .ZN(n_0_453));
   AND2_X1 i_0_0_173 (.A1(n_0_305), .A2(n_0_561), .ZN(n_0_454));
   AND2_X1 i_0_0_174 (.A1(n_0_306), .A2(n_0_561), .ZN(n_0_455));
   AND2_X1 i_0_0_175 (.A1(n_0_307), .A2(n_0_561), .ZN(n_0_456));
   AND2_X1 i_0_0_176 (.A1(n_0_308), .A2(n_0_561), .ZN(n_0_457));
   AND2_X1 i_0_0_177 (.A1(n_0_309), .A2(n_0_561), .ZN(n_0_487));
   AND2_X1 i_0_0_178 (.A1(n_0_310), .A2(n_0_561), .ZN(n_0_488));
   AND2_X1 i_0_0_179 (.A1(n_0_311), .A2(n_0_561), .ZN(n_0_489));
   AND2_X1 i_0_0_180 (.A1(n_0_312), .A2(n_0_561), .ZN(n_0_490));
   AND2_X1 i_0_0_181 (.A1(n_0_313), .A2(n_0_561), .ZN(n_0_491));
   AND2_X1 i_0_0_182 (.A1(n_0_314), .A2(n_0_561), .ZN(n_0_492));
   AND2_X1 i_0_0_183 (.A1(n_0_315), .A2(n_0_561), .ZN(n_0_493));
   AND2_X1 i_0_0_184 (.A1(n_0_316), .A2(n_0_561), .ZN(n_0_494));
   AND2_X1 i_0_0_185 (.A1(n_0_317), .A2(n_0_561), .ZN(n_0_495));
   AND2_X1 i_0_0_186 (.A1(n_0_318), .A2(n_0_561), .ZN(n_0_496));
   AND2_X1 i_0_0_187 (.A1(n_0_319), .A2(n_0_561), .ZN(n_0_497));
   AND2_X1 i_0_0_188 (.A1(n_0_320), .A2(n_0_561), .ZN(n_0_498));
   AND2_X1 i_0_0_189 (.A1(n_0_321), .A2(n_0_561), .ZN(n_0_499));
   AND2_X1 i_0_0_190 (.A1(n_0_322), .A2(n_0_561), .ZN(n_0_500));
   AND2_X1 i_0_0_191 (.A1(n_0_323), .A2(n_0_561), .ZN(n_0_501));
   AND2_X1 i_0_0_192 (.A1(n_0_324), .A2(n_0_561), .ZN(n_0_502));
   AND2_X1 i_0_0_193 (.A1(n_0_325), .A2(n_0_561), .ZN(n_0_503));
   OAI21_X1 i_0_0_194 (.A(n_0_0_73), .B1(n_0_0_370), .B2(n_0_0_208), .ZN(n_0_504));
   NOR3_X1 i_0_0_195 (.A1(n_0_0_275), .A2(reset), .A3(filterCounter[0]), 
      .ZN(n_0_0));
   AND2_X1 i_0_0_196 (.A1(n_0_230), .A2(n_0_0_83), .ZN(n_0_4));
   AND2_X1 i_0_0_197 (.A1(n_0_231), .A2(n_0_0_83), .ZN(n_0_10));
   AND2_X1 i_0_0_198 (.A1(n_0_232), .A2(n_0_0_83), .ZN(n_0_11));
   AND2_X1 i_0_0_199 (.A1(n_0_233), .A2(n_0_0_83), .ZN(n_0_12));
   AND2_X1 i_0_0_200 (.A1(n_0_235), .A2(n_0_0_83), .ZN(n_0_13));
   AND2_X1 i_0_0_201 (.A1(n_0_236), .A2(n_0_0_83), .ZN(n_0_17));
   AND2_X1 i_0_0_202 (.A1(n_0_237), .A2(n_0_0_83), .ZN(n_0_18));
   AND2_X1 i_0_0_203 (.A1(n_0_238), .A2(n_0_0_83), .ZN(n_0_19));
   AND2_X1 i_0_0_204 (.A1(n_0_239), .A2(n_0_0_83), .ZN(n_0_20));
   AND2_X1 i_0_0_205 (.A1(n_0_240), .A2(n_0_0_83), .ZN(n_0_21));
   AND2_X1 i_0_0_206 (.A1(n_0_241), .A2(n_0_0_83), .ZN(n_0_22));
   AND2_X1 i_0_0_207 (.A1(n_0_242), .A2(n_0_0_83), .ZN(n_0_24));
   AND2_X1 i_0_0_208 (.A1(n_0_243), .A2(n_0_0_83), .ZN(n_0_505));
   AND2_X1 i_0_0_209 (.A1(n_0_244), .A2(n_0_0_83), .ZN(n_0_506));
   AND2_X1 i_0_0_210 (.A1(n_0_245), .A2(n_0_0_83), .ZN(n_0_507));
   AND2_X1 i_0_0_211 (.A1(n_0_246), .A2(n_0_0_83), .ZN(n_0_508));
   AND2_X1 i_0_0_212 (.A1(n_0_247), .A2(n_0_0_83), .ZN(n_0_509));
   AND2_X1 i_0_0_213 (.A1(n_0_248), .A2(n_0_0_83), .ZN(n_0_511));
   AND2_X1 i_0_0_214 (.A1(n_0_249), .A2(n_0_0_83), .ZN(n_0_512));
   AND2_X1 i_0_0_215 (.A1(n_0_250), .A2(n_0_0_83), .ZN(n_0_513));
   AND2_X1 i_0_0_216 (.A1(n_0_251), .A2(n_0_0_83), .ZN(n_0_514));
   AND2_X1 i_0_0_217 (.A1(n_0_252), .A2(n_0_0_83), .ZN(n_0_515));
   AND2_X1 i_0_0_218 (.A1(n_0_253), .A2(n_0_0_83), .ZN(n_0_516));
   AND2_X1 i_0_0_219 (.A1(n_0_254), .A2(n_0_0_83), .ZN(n_0_517));
   AND2_X1 i_0_0_220 (.A1(n_0_255), .A2(n_0_0_83), .ZN(n_0_518));
   AND2_X1 i_0_0_221 (.A1(n_0_256), .A2(n_0_0_83), .ZN(n_0_519));
   AND2_X1 i_0_0_222 (.A1(n_0_257), .A2(n_0_0_83), .ZN(n_0_520));
   AND2_X1 i_0_0_223 (.A1(n_0_258), .A2(n_0_0_83), .ZN(n_0_521));
   AND2_X1 i_0_0_224 (.A1(n_0_259), .A2(n_0_0_83), .ZN(n_0_522));
   AND2_X1 i_0_0_225 (.A1(n_0_260), .A2(n_0_0_83), .ZN(n_0_523));
   AND2_X1 i_0_0_226 (.A1(n_0_261), .A2(n_0_0_83), .ZN(n_0_524));
   NOR2_X1 i_0_0_227 (.A1(n_0_0_275), .A2(reset), .ZN(n_0_0_83));
   NOR2_X1 i_0_0_228 (.A1(n_0_0_268), .A2(n_0_0_84), .ZN(n_0_557));
   NAND2_X1 i_0_0_229 (.A1(n_0_0_73), .A2(DMA_start), .ZN(n_0_0_84));
   OR2_X1 i_0_0_230 (.A1(n_0_0_347), .A2(n_0_553), .ZN(n_0_559));
   OAI21_X1 i_0_0_231 (.A(n_0_0_73), .B1(n_0_0_303), .B2(n_0_0_283), .ZN(n_0_553));
   OAI21_X1 i_0_0_232 (.A(n_0_0_73), .B1(n_0_0_435), .B2(n_0_0_432), .ZN(n_0_560));
   INV_X1 i_0_0_240 (.A(n_0_0_87), .ZN(n_0_36));
   AOI21_X1 i_0_0_241 (.A(reset), .B1(convState), .B2(n_0_0_88), .ZN(n_0_0_87));
   OR2_X1 i_0_0_242 (.A1(reset), .A2(n_0_0_88), .ZN(n_0_558));
   NOR3_X1 i_0_0_243 (.A1(n_0_0_275), .A2(n_0_0_208), .A3(n_0_0_389), .ZN(
      n_0_0_88));
   OAI21_X1 i_0_0_244 (.A(n_0_0_89), .B1(n_0_0_127), .B2(n_0_585), .ZN(n_0_38));
   AOI222_X1 i_0_0_245 (.A1(n_0_681), .A2(n_0_0_277), .B1(n_0_0_270), .B2(
      n_0_181), .C1(n_0_78), .C2(n_0_0_131), .ZN(n_0_0_89));
   AOI211_X1 i_0_0_246 (.A(n_0_0_91), .B(n_0_0_90), .C1(n_0_682), .C2(n_0_0_277), 
      .ZN(n_0_39));
   NOR2_X1 i_0_0_247 (.A1(n_0_0_130), .A2(n_0_79), .ZN(n_0_0_90));
   AOI221_X1 i_0_0_248 (.A(n_0_0_92), .B1(n_0_0_273), .B2(n_0_182), .C1(n_0_57), 
      .C2(n_0_0_134), .ZN(n_0_0_91));
   OAI211_X1 i_0_0_249 (.A(n_0_0_93), .B(n_0_0_431), .C1(n_0_0_454), .C2(
      n_0_0_110), .ZN(n_0_0_92));
   OAI21_X1 i_0_0_250 (.A(n_0_0_397), .B1(n_0_0_449), .B2(n_0_548), .ZN(n_0_0_93));
   OAI21_X1 i_0_0_251 (.A(n_0_0_94), .B1(n_0_0_95), .B2(n_0_0_96), .ZN(n_0_40));
   AOI22_X1 i_0_0_252 (.A1(n_0_0_31), .A2(n_0_0_277), .B1(n_0_0_131), .B2(n_0_80), 
      .ZN(n_0_0_94));
   OAI211_X1 i_0_0_253 (.A(n_0_0_431), .B(n_0_0_97), .C1(n_0_0_133), .C2(n_0_58), 
      .ZN(n_0_0_95));
   NOR2_X1 i_0_0_254 (.A1(n_0_0_272), .A2(n_0_183), .ZN(n_0_0_96));
   OAI21_X1 i_0_0_255 (.A(n_0_0_397), .B1(n_0_0_424), .B2(n_0_570), .ZN(n_0_0_97));
   NOR2_X1 i_0_0_256 (.A1(n_0_0_98), .A2(n_0_0_100), .ZN(n_0_41));
   AOI221_X1 i_0_0_257 (.A(n_0_0_99), .B1(n_0_0_273), .B2(n_0_200), .C1(n_0_59), 
      .C2(n_0_0_134), .ZN(n_0_0_98));
   OAI21_X1 i_0_0_258 (.A(n_0_0_431), .B1(n_0_0_381), .B2(n_0_0_110), .ZN(
      n_0_0_99));
   OAI22_X1 i_0_0_259 (.A1(n_0_0_32), .A2(n_0_0_276), .B1(n_0_0_130), .B2(n_0_81), 
      .ZN(n_0_0_100));
   AOI211_X1 i_0_0_260 (.A(n_0_0_104), .B(n_0_0_101), .C1(n_0_0_102), .C2(
      n_0_568), .ZN(n_0_42));
   OAI22_X1 i_0_0_261 (.A1(n_0_0_127), .A2(n_0_60), .B1(n_0_0_269), .B2(n_0_201), 
      .ZN(n_0_0_101));
   XNOR2_X1 i_0_0_262 (.A(n_0_0_86), .B(n_0_0_103), .ZN(n_0_0_102));
   NOR2_X1 i_0_0_263 (.A1(n_0_0_65), .A2(convResetState[0]), .ZN(n_0_0_103));
   OAI22_X1 i_0_0_264 (.A1(n_0_0_33), .A2(n_0_0_276), .B1(n_0_0_130), .B2(n_0_82), 
      .ZN(n_0_0_104));
   NOR2_X1 i_0_0_265 (.A1(n_0_0_106), .A2(n_0_0_105), .ZN(n_0_43));
   OAI22_X1 i_0_0_266 (.A1(n_0_0_34), .A2(n_0_0_276), .B1(n_0_0_130), .B2(n_0_83), 
      .ZN(n_0_0_105));
   AOI221_X1 i_0_0_267 (.A(n_0_0_109), .B1(n_0_0_273), .B2(n_0_202), .C1(n_0_61), 
      .C2(n_0_0_134), .ZN(n_0_0_106));
   NOR2_X1 i_0_0_268 (.A1(n_0_0_108), .A2(n_0_0_107), .ZN(n_0_44));
   OAI22_X1 i_0_0_269 (.A1(n_0_0_35), .A2(n_0_0_276), .B1(n_0_0_130), .B2(n_0_84), 
      .ZN(n_0_0_107));
   AOI221_X1 i_0_0_270 (.A(n_0_0_109), .B1(n_0_0_273), .B2(n_0_203), .C1(n_0_62), 
      .C2(n_0_0_134), .ZN(n_0_0_108));
   OAI221_X1 i_0_0_271 (.A(n_0_0_431), .B1(n_0_0_110), .B2(layerCounter[2]), 
      .C1(n_0_0_428), .C2(n_0_0_448), .ZN(n_0_0_109));
   NAND2_X1 i_0_0_272 (.A1(n_0_0_72), .A2(convResetState[0]), .ZN(n_0_0_110));
   NOR3_X1 i_0_0_273 (.A1(n_0_0_114), .A2(n_0_0_113), .A3(n_0_0_111), .ZN(n_0_45));
   OAI221_X1 i_0_0_274 (.A(n_0_0_112), .B1(n_0_0_276), .B2(n_0_0_36), .C1(n_0_85), 
      .C2(n_0_0_130), .ZN(n_0_0_111));
   OAI211_X1 i_0_0_275 (.A(n_0_568), .B(n_0_0_462), .C1(convResetState[0]), 
      .C2(n_0_0_456), .ZN(n_0_0_112));
   NOR2_X1 i_0_0_276 (.A1(n_0_0_269), .A2(n_0_204), .ZN(n_0_0_113));
   NOR2_X1 i_0_0_277 (.A1(n_0_0_127), .A2(n_0_63), .ZN(n_0_0_114));
   NAND2_X1 i_0_0_278 (.A1(n_0_0_115), .A2(n_0_0_117), .ZN(n_0_46));
   OAI221_X1 i_0_0_279 (.A(n_0_0_116), .B1(n_0_0_133), .B2(n_0_64), .C1(
      n_0_0_272), .C2(n_0_205), .ZN(n_0_0_115));
   AOI21_X1 i_0_0_280 (.A(n_0_0_430), .B1(n_0_0_397), .B2(n_0_0_462), .ZN(
      n_0_0_116));
   AOI22_X1 i_0_0_281 (.A1(n_0_0_37), .A2(n_0_0_277), .B1(n_0_0_131), .B2(n_0_86), 
      .ZN(n_0_0_117));
   OAI21_X1 i_0_0_282 (.A(n_0_0_118), .B1(n_0_0_127), .B2(n_0_0_475), .ZN(n_0_47));
   AOI222_X1 i_0_0_283 (.A1(n_0_0_38), .A2(n_0_0_277), .B1(n_0_0_270), .B2(
      n_0_206), .C1(n_0_87), .C2(n_0_0_131), .ZN(n_0_0_118));
   NOR2_X1 i_0_0_284 (.A1(n_0_0_120), .A2(n_0_0_119), .ZN(n_0_48));
   OAI22_X1 i_0_0_285 (.A1(n_0_0_127), .A2(n_0_66), .B1(n_0_0_269), .B2(n_0_207), 
      .ZN(n_0_0_119));
   AOI221_X1 i_0_0_286 (.A(n_0_0_135), .B1(n_0_0_131), .B2(n_0_88), .C1(n_0_0_39), 
      .C2(n_0_0_277), .ZN(n_0_0_120));
   AOI21_X1 i_0_0_287 (.A(n_0_0_121), .B1(n_0_0_122), .B2(n_0_0_123), .ZN(n_0_49));
   OAI22_X1 i_0_0_288 (.A1(n_0_0_40), .A2(n_0_0_276), .B1(n_0_0_130), .B2(n_0_89), 
      .ZN(n_0_0_121));
   AOI221_X1 i_0_0_289 (.A(n_0_0_430), .B1(n_0_0_397), .B2(n_0_0_449), .C1(
      n_0_0_134), .C2(n_0_67), .ZN(n_0_0_122));
   NAND2_X1 i_0_0_290 (.A1(n_0_208), .A2(n_0_0_273), .ZN(n_0_0_123));
   OAI21_X1 i_0_0_291 (.A(n_0_0_124), .B1(n_0_0_127), .B2(n_0_0_67), .ZN(n_0_50));
   AOI222_X1 i_0_0_292 (.A1(n_0_0_41), .A2(n_0_0_277), .B1(n_0_0_270), .B2(
      n_0_209), .C1(n_0_90), .C2(n_0_0_131), .ZN(n_0_0_124));
   OAI21_X1 i_0_0_293 (.A(n_0_0_125), .B1(n_0_0_127), .B2(n_0_0_68), .ZN(n_0_51));
   AOI222_X1 i_0_0_294 (.A1(n_0_0_42), .A2(n_0_0_277), .B1(n_0_0_270), .B2(
      n_0_210), .C1(n_0_91), .C2(n_0_0_131), .ZN(n_0_0_125));
   NOR2_X1 i_0_0_295 (.A1(n_0_0_128), .A2(n_0_0_126), .ZN(n_0_52));
   OAI22_X1 i_0_0_296 (.A1(n_0_0_127), .A2(n_0_70), .B1(n_0_0_269), .B2(n_0_211), 
      .ZN(n_0_0_126));
   NAND2_X1 i_0_0_297 (.A1(n_0_0_275), .A2(n_0_0_271), .ZN(n_0_0_127));
   AOI221_X1 i_0_0_298 (.A(n_0_0_135), .B1(n_0_0_131), .B2(n_0_92), .C1(n_0_0_43), 
      .C2(n_0_0_277), .ZN(n_0_0_128));
   NAND2_X1 i_0_0_299 (.A1(n_0_0_132), .A2(n_0_0_129), .ZN(n_0_53));
   AOI22_X1 i_0_0_300 (.A1(n_0_0_277), .A2(n_0_0_171), .B1(n_0_0_131), .B2(
      n_0_93), .ZN(n_0_0_129));
   NAND2_X1 i_0_0_301 (.A1(n_0_0_430), .A2(n_0_0_278), .ZN(n_0_0_130));
   NOR2_X1 i_0_0_302 (.A1(n_0_0_431), .A2(n_0_0_429), .ZN(n_0_0_131));
   OAI221_X1 i_0_0_303 (.A(n_0_0_135), .B1(n_0_0_133), .B2(n_0_71), .C1(
      n_0_0_272), .C2(n_0_212), .ZN(n_0_0_132));
   NAND2_X1 i_0_0_304 (.A1(n_0_0_275), .A2(convResetState[1]), .ZN(n_0_0_133));
   NOR2_X1 i_0_0_305 (.A1(n_0_0_274), .A2(n_0_0_72), .ZN(n_0_0_134));
   NOR2_X1 i_0_0_306 (.A1(n_0_0_430), .A2(n_0_0_397), .ZN(n_0_0_135));
   NOR2_X1 i_0_0_307 (.A1(n_0_0_389), .A2(n_0_0_214), .ZN(n_0_561));
   OAI21_X1 i_0_0_308 (.A(n_0_0_73), .B1(n_0_0_136), .B2(n_0_0_208), .ZN(n_0_562));
   NOR2_X1 i_0_0_309 (.A1(n_0_0_389), .A2(n_0_0_469), .ZN(n_0_0_136));
   NAND2_X1 i_0_0_310 (.A1(n_0_0_138), .A2(n_0_0_137), .ZN(n_0_54));
   AOI222_X1 i_0_0_311 (.A1(n_0_0_175), .A2(n_0_697), .B1(n_0_0_264), .B2(
      n_0_181), .C1(n_0_0_173), .C2(n_0_165), .ZN(n_0_0_137));
   AOI22_X1 i_0_0_312 (.A1(n_0_111), .A2(n_0_0_172), .B1(n_0_0_177), .B2(n_0_681), 
      .ZN(n_0_0_138));
   NAND2_X1 i_0_0_313 (.A1(n_0_0_140), .A2(n_0_0_139), .ZN(n_0_55));
   AOI22_X1 i_0_0_314 (.A1(n_0_0_175), .A2(n_0_698), .B1(n_0_0_264), .B2(n_0_182), 
      .ZN(n_0_0_139));
   AOI221_X1 i_0_0_315 (.A(n_0_0_141), .B1(n_0_0_173), .B2(n_0_166), .C1(n_0_112), 
      .C2(n_0_0_172), .ZN(n_0_0_140));
   MUX2_X1 i_0_0_316 (.A(n_0_0_260), .B(n_0_0_176), .S(n_0_682), .Z(n_0_0_141));
   NAND2_X1 i_0_0_317 (.A1(n_0_0_143), .A2(n_0_0_142), .ZN(n_0_276));
   AOI222_X1 i_0_0_318 (.A1(n_0_0_175), .A2(n_0_699), .B1(n_0_0_264), .B2(
      n_0_183), .C1(n_0_0_173), .C2(n_0_167), .ZN(n_0_0_142));
   AOI222_X1 i_0_0_319 (.A1(n_0_0_31), .A2(n_0_0_260), .B1(n_0_0_172), .B2(
      n_0_113), .C1(n_0_683), .C2(n_0_0_176), .ZN(n_0_0_143));
   NAND2_X1 i_0_0_320 (.A1(n_0_0_145), .A2(n_0_0_144), .ZN(n_0_277));
   AOI222_X1 i_0_0_321 (.A1(n_0_0_175), .A2(n_0_1), .B1(n_0_0_264), .B2(n_0_200), 
      .C1(n_0_0_173), .C2(n_0_168), .ZN(n_0_0_144));
   AOI222_X1 i_0_0_322 (.A1(n_0_0_32), .A2(n_0_0_260), .B1(n_0_0_172), .B2(
      n_0_114), .C1(n_0_684), .C2(n_0_0_176), .ZN(n_0_0_145));
   NAND2_X1 i_0_0_323 (.A1(n_0_0_147), .A2(n_0_0_146), .ZN(n_0_278));
   AOI222_X1 i_0_0_324 (.A1(n_0_0_175), .A2(n_0_3), .B1(n_0_0_264), .B2(n_0_201), 
      .C1(n_0_0_173), .C2(n_0_169), .ZN(n_0_0_146));
   AOI222_X1 i_0_0_325 (.A1(n_0_0_33), .A2(n_0_0_260), .B1(n_0_0_172), .B2(
      n_0_115), .C1(n_0_685), .C2(n_0_0_176), .ZN(n_0_0_147));
   NAND2_X1 i_0_0_326 (.A1(n_0_0_149), .A2(n_0_0_148), .ZN(n_0_280));
   AOI222_X1 i_0_0_327 (.A1(n_0_0_175), .A2(n_0_25), .B1(n_0_0_264), .B2(n_0_202), 
      .C1(n_0_0_173), .C2(n_0_170), .ZN(n_0_0_148));
   AOI222_X1 i_0_0_328 (.A1(n_0_0_34), .A2(n_0_0_260), .B1(n_0_0_172), .B2(
      n_0_116), .C1(n_0_686), .C2(n_0_0_176), .ZN(n_0_0_149));
   NAND2_X1 i_0_0_329 (.A1(n_0_0_151), .A2(n_0_0_150), .ZN(n_0_281));
   AOI222_X1 i_0_0_330 (.A1(n_0_0_175), .A2(n_0_30), .B1(n_0_0_264), .B2(n_0_203), 
      .C1(n_0_0_173), .C2(n_0_171), .ZN(n_0_0_150));
   AOI222_X1 i_0_0_331 (.A1(n_0_0_35), .A2(n_0_0_260), .B1(n_0_0_172), .B2(
      n_0_117), .C1(n_0_687), .C2(n_0_0_176), .ZN(n_0_0_151));
   NAND2_X1 i_0_0_332 (.A1(n_0_0_153), .A2(n_0_0_152), .ZN(n_0_282));
   AOI222_X1 i_0_0_333 (.A1(n_0_0_175), .A2(n_0_31), .B1(n_0_0_264), .B2(n_0_204), 
      .C1(n_0_0_173), .C2(n_0_172), .ZN(n_0_0_152));
   AOI222_X1 i_0_0_334 (.A1(n_0_0_36), .A2(n_0_0_260), .B1(n_0_0_172), .B2(
      n_0_118), .C1(n_0_688), .C2(n_0_0_176), .ZN(n_0_0_153));
   NAND2_X1 i_0_0_335 (.A1(n_0_0_155), .A2(n_0_0_154), .ZN(n_0_525));
   AOI222_X1 i_0_0_336 (.A1(n_0_0_175), .A2(n_0_32), .B1(n_0_0_264), .B2(n_0_205), 
      .C1(n_0_0_173), .C2(n_0_173), .ZN(n_0_0_154));
   AOI222_X1 i_0_0_337 (.A1(n_0_0_37), .A2(n_0_0_260), .B1(n_0_0_172), .B2(
      n_0_119), .C1(n_0_689), .C2(n_0_0_176), .ZN(n_0_0_155));
   NAND2_X1 i_0_0_338 (.A1(n_0_0_157), .A2(n_0_0_156), .ZN(n_0_526));
   AOI222_X1 i_0_0_339 (.A1(n_0_0_175), .A2(n_0_34), .B1(n_0_0_264), .B2(n_0_206), 
      .C1(n_0_0_173), .C2(n_0_174), .ZN(n_0_0_156));
   AOI222_X1 i_0_0_340 (.A1(n_0_0_38), .A2(n_0_0_260), .B1(n_0_0_172), .B2(
      n_0_130), .C1(n_0_690), .C2(n_0_0_176), .ZN(n_0_0_157));
   NAND2_X1 i_0_0_341 (.A1(n_0_0_159), .A2(n_0_0_158), .ZN(n_0_527));
   AOI222_X1 i_0_0_342 (.A1(n_0_0_175), .A2(n_0_533), .B1(n_0_0_264), .B2(
      n_0_207), .C1(n_0_0_173), .C2(n_0_175), .ZN(n_0_0_158));
   AOI222_X1 i_0_0_343 (.A1(n_0_0_39), .A2(n_0_0_260), .B1(n_0_0_172), .B2(
      n_0_131), .C1(n_0_691), .C2(n_0_0_176), .ZN(n_0_0_159));
   NAND2_X1 i_0_0_344 (.A1(n_0_0_161), .A2(n_0_0_160), .ZN(n_0_528));
   AOI222_X1 i_0_0_345 (.A1(n_0_0_175), .A2(n_0_534), .B1(n_0_0_264), .B2(
      n_0_208), .C1(n_0_0_173), .C2(n_0_176), .ZN(n_0_0_160));
   AOI222_X1 i_0_0_346 (.A1(n_0_0_40), .A2(n_0_0_260), .B1(n_0_0_172), .B2(
      n_0_132), .C1(n_0_692), .C2(n_0_0_176), .ZN(n_0_0_161));
   NAND2_X1 i_0_0_347 (.A1(n_0_0_163), .A2(n_0_0_162), .ZN(n_0_529));
   AOI222_X1 i_0_0_348 (.A1(n_0_0_175), .A2(n_0_535), .B1(n_0_0_264), .B2(
      n_0_209), .C1(n_0_0_173), .C2(n_0_177), .ZN(n_0_0_162));
   AOI222_X1 i_0_0_349 (.A1(n_0_0_41), .A2(n_0_0_260), .B1(n_0_0_172), .B2(
      n_0_133), .C1(n_0_693), .C2(n_0_0_176), .ZN(n_0_0_163));
   NAND2_X1 i_0_0_350 (.A1(n_0_0_165), .A2(n_0_0_164), .ZN(n_0_530));
   AOI222_X1 i_0_0_351 (.A1(n_0_0_175), .A2(n_0_536), .B1(n_0_0_264), .B2(
      n_0_210), .C1(n_0_0_173), .C2(n_0_178), .ZN(n_0_0_164));
   AOI222_X1 i_0_0_352 (.A1(n_0_0_42), .A2(n_0_0_260), .B1(n_0_0_172), .B2(
      n_0_134), .C1(n_0_694), .C2(n_0_0_176), .ZN(n_0_0_165));
   NAND2_X1 i_0_0_353 (.A1(n_0_0_167), .A2(n_0_0_166), .ZN(n_0_531));
   AOI222_X1 i_0_0_354 (.A1(n_0_0_175), .A2(n_0_537), .B1(n_0_0_264), .B2(
      n_0_211), .C1(n_0_0_173), .C2(n_0_179), .ZN(n_0_0_166));
   AOI222_X1 i_0_0_355 (.A1(n_0_0_43), .A2(n_0_0_260), .B1(n_0_0_172), .B2(
      n_0_135), .C1(n_0_695), .C2(n_0_0_176), .ZN(n_0_0_167));
   NAND2_X1 i_0_0_356 (.A1(n_0_0_174), .A2(n_0_0_168), .ZN(n_0_532));
   AOI221_X1 i_0_0_357 (.A(n_0_0_169), .B1(n_0_0_176), .B2(n_0_696), .C1(n_0_180), 
      .C2(n_0_0_173), .ZN(n_0_0_168));
   INV_X1 i_0_0_358 (.A(n_0_0_170), .ZN(n_0_0_169));
   AOI22_X1 i_0_0_359 (.A1(n_0_136), .A2(n_0_0_172), .B1(n_0_0_171), .B2(
      n_0_0_260), .ZN(n_0_0_170));
   XOR2_X1 i_0_0_360 (.A(n_0_0_13), .B(n_0_696), .Z(n_0_0_171));
   NOR2_X1 i_0_0_361 (.A1(n_0_0_282), .A2(n_0_0_262), .ZN(n_0_0_172));
   AND2_X1 i_0_0_362 (.A1(n_0_0_431), .A2(n_0_0_204), .ZN(n_0_0_173));
   AOI22_X1 i_0_0_363 (.A1(n_0_0_175), .A2(n_0_538), .B1(n_0_0_264), .B2(n_0_212), 
      .ZN(n_0_0_174));
   NOR3_X1 i_0_0_364 (.A1(n_0_0_265), .A2(n_0_0_204), .A3(n_0_0_430), .ZN(
      n_0_0_175));
   OAI21_X1 i_0_0_365 (.A(n_0_0_179), .B1(n_0_0_178), .B2(n_0_0_261), .ZN(
      n_0_0_176));
   NAND2_X1 i_0_0_366 (.A1(n_0_0_179), .A2(n_0_0_178), .ZN(n_0_0_177));
   NAND2_X1 i_0_0_367 (.A1(n_0_0_282), .A2(layerCounter[0]), .ZN(n_0_0_178));
   NAND2_X1 i_0_0_368 (.A1(n_0_0_430), .A2(n_0_0_263), .ZN(n_0_0_179));
   OAI21_X1 i_0_0_369 (.A(n_0_0_180), .B1(n_0_0_452), .B2(convReset), .ZN(
      n_0_697));
   NAND2_X1 i_0_0_370 (.A1(convReset), .A2(readAdress[0]), .ZN(n_0_0_180));
   OAI21_X1 i_0_0_371 (.A(n_0_0_181), .B1(n_0_0_452), .B2(convReset), .ZN(
      n_0_698));
   NAND2_X1 i_0_0_372 (.A1(convReset), .A2(readAdress[1]), .ZN(n_0_0_181));
   OAI21_X1 i_0_0_373 (.A(n_0_0_182), .B1(n_0_539), .B2(convReset), .ZN(n_0_699));
   NAND2_X1 i_0_0_374 (.A1(convReset), .A2(readAdress[2]), .ZN(n_0_0_182));
   MUX2_X1 i_0_0_375 (.A(n_0_0_44), .B(readAdress[3]), .S(convReset), .Z(n_0_1));
   MUX2_X1 i_0_0_376 (.A(n_0_0_45), .B(readAdress[4]), .S(convReset), .Z(n_0_3));
   MUX2_X1 i_0_0_377 (.A(n_0_0_46), .B(readAdress[5]), .S(convReset), .Z(n_0_25));
   MUX2_X1 i_0_0_378 (.A(n_0_0_47), .B(readAdress[6]), .S(convReset), .Z(n_0_30));
   MUX2_X1 i_0_0_379 (.A(n_0_0_48), .B(readAdress[7]), .S(convReset), .Z(n_0_31));
   MUX2_X1 i_0_0_380 (.A(n_0_0_49), .B(readAdress[8]), .S(convReset), .Z(n_0_32));
   MUX2_X1 i_0_0_381 (.A(n_0_0_50), .B(readAdress[9]), .S(convReset), .Z(n_0_34));
   MUX2_X1 i_0_0_382 (.A(n_0_0_51), .B(readAdress[10]), .S(convReset), .Z(
      n_0_533));
   MUX2_X1 i_0_0_383 (.A(n_0_0_52), .B(readAdress[11]), .S(convReset), .Z(
      n_0_534));
   MUX2_X1 i_0_0_384 (.A(n_0_0_53), .B(readAdress[12]), .S(convReset), .Z(
      n_0_535));
   MUX2_X1 i_0_0_385 (.A(n_0_0_54), .B(readAdress[13]), .S(convReset), .Z(
      n_0_536));
   OAI21_X1 i_0_0_386 (.A(n_0_0_183), .B1(n_0_0_467), .B2(n_0_0_469), .ZN(
      n_0_537));
   OAI21_X1 i_0_0_387 (.A(n_0_0_183), .B1(n_0_0_468), .B2(n_0_0_469), .ZN(
      n_0_538));
   NAND2_X1 i_0_0_388 (.A1(n_0_0_469), .A2(n_0_0_184), .ZN(n_0_0_183));
   XNOR2_X1 i_0_0_389 (.A(n_0_0_24), .B(n_0_0_58), .ZN(n_0_0_184));
   MUX2_X1 i_0_0_390 (.A(n_0_0_204), .B(n_0_0_203), .S(n_0_649), .Z(n_0_665));
   OAI21_X1 i_0_0_391 (.A(n_0_0_186), .B1(n_0_0_185), .B2(n_0_0_204), .ZN(
      n_0_666));
   NAND2_X1 i_0_0_392 (.A1(n_0_0_371), .A2(n_0_650), .ZN(n_0_0_185));
   NAND2_X1 i_0_0_393 (.A1(n_0_95), .A2(n_0_0_204), .ZN(n_0_0_186));
   INV_X1 i_0_0_394 (.A(n_0_0_187), .ZN(n_0_667));
   AOI22_X1 i_0_0_395 (.A1(n_0_0_203), .A2(n_0_651), .B1(n_0_96), .B2(n_0_0_204), 
      .ZN(n_0_0_187));
   NAND2_X1 i_0_0_396 (.A1(n_0_0_189), .A2(n_0_0_188), .ZN(n_0_668));
   NAND2_X1 i_0_0_397 (.A1(n_0_652), .A2(n_0_0_203), .ZN(n_0_0_188));
   NAND2_X1 i_0_0_398 (.A1(n_0_97), .A2(n_0_0_204), .ZN(n_0_0_189));
   INV_X1 i_0_0_399 (.A(n_0_0_190), .ZN(n_0_669));
   AOI22_X1 i_0_0_400 (.A1(n_0_98), .A2(n_0_0_204), .B1(n_0_0_203), .B2(n_0_653), 
      .ZN(n_0_0_190));
   INV_X1 i_0_0_401 (.A(n_0_0_191), .ZN(n_0_670));
   AOI22_X1 i_0_0_402 (.A1(n_0_99), .A2(n_0_0_204), .B1(n_0_0_203), .B2(n_0_654), 
      .ZN(n_0_0_191));
   INV_X1 i_0_0_403 (.A(n_0_0_192), .ZN(n_0_671));
   AOI22_X1 i_0_0_404 (.A1(n_0_100), .A2(n_0_0_204), .B1(n_0_0_203), .B2(n_0_655), 
      .ZN(n_0_0_192));
   INV_X1 i_0_0_405 (.A(n_0_0_193), .ZN(n_0_672));
   AOI22_X1 i_0_0_406 (.A1(n_0_0_203), .A2(n_0_656), .B1(n_0_101), .B2(n_0_0_204), 
      .ZN(n_0_0_193));
   INV_X1 i_0_0_407 (.A(n_0_0_194), .ZN(n_0_673));
   AOI22_X1 i_0_0_408 (.A1(n_0_0_203), .A2(n_0_657), .B1(n_0_102), .B2(n_0_0_204), 
      .ZN(n_0_0_194));
   INV_X1 i_0_0_409 (.A(n_0_0_195), .ZN(n_0_674));
   AOI22_X1 i_0_0_410 (.A1(n_0_0_203), .A2(n_0_658), .B1(n_0_103), .B2(n_0_0_204), 
      .ZN(n_0_0_195));
   INV_X1 i_0_0_411 (.A(n_0_0_196), .ZN(n_0_675));
   AOI22_X1 i_0_0_412 (.A1(n_0_0_203), .A2(n_0_659), .B1(n_0_104), .B2(n_0_0_204), 
      .ZN(n_0_0_196));
   INV_X1 i_0_0_413 (.A(n_0_0_197), .ZN(n_0_676));
   AOI22_X1 i_0_0_414 (.A1(n_0_105), .A2(n_0_0_204), .B1(n_0_0_203), .B2(n_0_660), 
      .ZN(n_0_0_197));
   INV_X1 i_0_0_415 (.A(n_0_0_198), .ZN(n_0_677));
   AOI22_X1 i_0_0_416 (.A1(n_0_0_203), .A2(n_0_661), .B1(n_0_106), .B2(n_0_0_204), 
      .ZN(n_0_0_198));
   NAND2_X1 i_0_0_417 (.A1(n_0_0_200), .A2(n_0_0_199), .ZN(n_0_678));
   NAND2_X1 i_0_0_418 (.A1(n_0_662), .A2(n_0_0_203), .ZN(n_0_0_199));
   NAND2_X1 i_0_0_419 (.A1(n_0_107), .A2(n_0_0_204), .ZN(n_0_0_200));
   INV_X1 i_0_0_420 (.A(n_0_0_201), .ZN(n_0_679));
   AOI22_X1 i_0_0_421 (.A1(n_0_0_203), .A2(n_0_663), .B1(n_0_108), .B2(n_0_0_204), 
      .ZN(n_0_0_201));
   INV_X1 i_0_0_422 (.A(n_0_0_202), .ZN(n_0_680));
   AOI22_X1 i_0_0_423 (.A1(n_0_0_203), .A2(n_0_664), .B1(n_0_109), .B2(n_0_0_204), 
      .ZN(n_0_0_202));
   NOR2_X1 i_0_0_424 (.A1(n_0_0_372), .A2(n_0_0_204), .ZN(n_0_0_203));
   AND3_X1 i_0_0_425 (.A1(DMA_start), .A2(n_0_0_369), .A3(n_0_0_349), .ZN(
      n_0_0_204));
   AND2_X1 i_0_0_426 (.A1(baseReadAdress[0]), .A2(convReset), .ZN(n_0_649));
   AND2_X1 i_0_0_427 (.A1(baseReadAdress[1]), .A2(convReset), .ZN(n_0_650));
   OR2_X1 i_0_0_428 (.A1(n_0_0_469), .A2(baseReadAdress[2]), .ZN(n_0_651));
   MUX2_X1 i_0_0_429 (.A(baseReadAdress[3]), .B(n_0_0_61), .S(n_0_0_469), 
      .Z(n_0_652));
   MUX2_X1 i_0_0_430 (.A(baseReadAdress[4]), .B(n_0_0_28), .S(n_0_0_469), 
      .Z(n_0_653));
   MUX2_X1 i_0_0_431 (.A(baseReadAdress[5]), .B(n_0_0_29), .S(n_0_0_469), 
      .Z(n_0_654));
   MUX2_X1 i_0_0_432 (.A(baseReadAdress[6]), .B(n_0_0_30), .S(n_0_0_469), 
      .Z(n_0_655));
   MUX2_X1 i_0_0_433 (.A(baseReadAdress[7]), .B(n_0_0_55), .S(n_0_0_469), 
      .Z(n_0_656));
   OAI21_X1 i_0_0_434 (.A(n_0_0_205), .B1(n_0_0_462), .B2(convReset), .ZN(
      n_0_657));
   NAND2_X1 i_0_0_435 (.A1(baseReadAdress[8]), .A2(convReset), .ZN(n_0_0_205));
   MUX2_X1 i_0_0_436 (.A(baseReadAdress[9]), .B(n_0_0_56), .S(n_0_0_469), 
      .Z(n_0_658));
   MUX2_X1 i_0_0_437 (.A(baseReadAdress[10]), .B(n_0_0_57), .S(n_0_0_469), 
      .Z(n_0_659));
   AOI21_X1 i_0_0_438 (.A(n_0_0_206), .B1(n_0_0_58), .B2(n_0_0_469), .ZN(n_0_660));
   NOR2_X1 i_0_0_439 (.A1(n_0_0_469), .A2(baseReadAdress[11]), .ZN(n_0_0_206));
   OAI21_X1 i_0_0_440 (.A(n_0_0_207), .B1(n_0_0_455), .B2(convReset), .ZN(
      n_0_661));
   NAND2_X1 i_0_0_441 (.A1(baseReadAdress[12]), .A2(convReset), .ZN(n_0_0_207));
   MUX2_X1 i_0_0_442 (.A(baseReadAdress[13]), .B(n_0_0_61), .S(n_0_0_469), 
      .Z(n_0_662));
   OR2_X1 i_0_0_443 (.A1(n_0_0_469), .A2(baseReadAdress[14]), .ZN(n_0_663));
   OR2_X1 i_0_0_444 (.A1(n_0_0_469), .A2(baseReadAdress[15]), .ZN(n_0_664));
   NOR2_X1 i_0_0_445 (.A1(n_0_0_208), .A2(reset), .ZN(n_0_638));
   NAND3_X1 i_0_0_446 (.A1(n_0_0_371), .A2(n_0_0_425), .A3(convResetState[1]), 
      .ZN(n_0_0_208));
   AOI21_X1 i_0_0_447 (.A(n_0_0_210), .B1(n_0_563), .B2(poolingReset), .ZN(
      n_0_564));
   INV_X1 i_0_0_448 (.A(n_0_563), .ZN(n_0_0_209));
   NOR2_X1 i_0_0_449 (.A1(reset), .A2(n_0_0_307), .ZN(n_0_563));
   AOI21_X1 i_0_0_450 (.A(reset), .B1(n_0_0_427), .B2(layerCounter[0]), .ZN(
      n_0_0_210));
   AOI211_X1 i_0_0_451 (.A(reset), .B(n_0_0_426), .C1(n_0_0_211), .C2(n_0_0_76), 
      .ZN(n_0_635));
   NAND2_X1 i_0_0_452 (.A1(n_0_0_371), .A2(convResetState[1]), .ZN(n_0_0_211));
   AOI21_X1 i_0_0_453 (.A(reset), .B1(n_0_0_372), .B2(n_0_0_271), .ZN(n_0_565));
   OAI21_X1 i_0_0_454 (.A(n_0_0_212), .B1(n_0_0_426), .B2(writeReset), .ZN(
      n_0_566));
   OR2_X1 i_0_0_455 (.A1(n_0_0_215), .A2(n_0_0_213), .ZN(n_0_0_212));
   AOI21_X1 i_0_0_456 (.A(reset), .B1(convResetState[1]), .B2(n_0_0_425), 
      .ZN(n_0_0_213));
   INV_X1 i_0_0_457 (.A(n_0_0_215), .ZN(n_0_0_214));
   NOR2_X1 i_0_0_458 (.A1(reset), .A2(n_0_0_372), .ZN(n_0_0_215));
   INV_X1 i_0_0_459 (.A(n_0_0_216), .ZN(n_0_617));
   MUX2_X1 i_0_0_460 (.A(n_0_0_240), .B(n_0_0_217), .S(n_0_0_247), .Z(n_0_0_216));
   AOI211_X1 i_0_0_461 (.A(n_0_0_239), .B(n_0_0_237), .C1(n_0_0_238), .C2(
      poolingReset), .ZN(n_0_0_217));
   OAI21_X1 i_0_0_462 (.A(n_0_0_218), .B1(n_0_0_240), .B2(n_0_0_248), .ZN(
      n_0_618));
   AOI221_X1 i_0_0_463 (.A(n_0_0_239), .B1(n_0_0_238), .B2(n_0_79), .C1(
      n_0_0_237), .C2(n_0_57), .ZN(n_0_0_218));
   NAND2_X1 i_0_0_464 (.A1(n_0_0_219), .A2(n_0_0_220), .ZN(n_0_619));
   AOI222_X1 i_0_0_465 (.A1(n_0_603), .A2(n_0_0_243), .B1(n_0_0_238), .B2(n_0_80), 
      .C1(n_0_58), .C2(n_0_0_237), .ZN(n_0_0_219));
   NAND2_X1 i_0_0_466 (.A1(n_0_587), .A2(n_0_0_241), .ZN(n_0_0_220));
   OAI21_X1 i_0_0_467 (.A(n_0_0_221), .B1(n_0_0_236), .B2(n_0_0_470), .ZN(
      n_0_620));
   AOI222_X1 i_0_0_468 (.A1(n_0_604), .A2(n_0_0_243), .B1(n_0_0_241), .B2(
      n_0_588), .C1(n_0_81), .C2(n_0_0_238), .ZN(n_0_0_221));
   OAI21_X1 i_0_0_469 (.A(n_0_0_222), .B1(n_0_0_236), .B2(n_0_0_471), .ZN(
      n_0_621));
   AOI222_X1 i_0_0_470 (.A1(n_0_0_241), .A2(n_0_589), .B1(n_0_82), .B2(n_0_0_238), 
      .C1(n_0_0_243), .C2(n_0_605), .ZN(n_0_0_222));
   OAI21_X1 i_0_0_471 (.A(n_0_0_223), .B1(n_0_0_236), .B2(n_0_0_472), .ZN(
      n_0_622));
   AOI222_X1 i_0_0_472 (.A1(n_0_0_241), .A2(n_0_590), .B1(n_0_83), .B2(n_0_0_238), 
      .C1(n_0_0_243), .C2(n_0_606), .ZN(n_0_0_223));
   OAI21_X1 i_0_0_473 (.A(n_0_0_224), .B1(n_0_0_236), .B2(n_0_0_473), .ZN(
      n_0_623));
   AOI222_X1 i_0_0_474 (.A1(n_0_607), .A2(n_0_0_243), .B1(n_0_0_241), .B2(
      n_0_591), .C1(n_0_84), .C2(n_0_0_238), .ZN(n_0_0_224));
   NAND2_X1 i_0_0_475 (.A1(n_0_0_225), .A2(n_0_0_226), .ZN(n_0_624));
   AOI222_X1 i_0_0_476 (.A1(n_0_85), .A2(n_0_0_238), .B1(n_0_0_237), .B2(n_0_63), 
      .C1(n_0_0_243), .C2(n_0_608), .ZN(n_0_0_225));
   NAND2_X1 i_0_0_477 (.A1(n_0_0_241), .A2(n_0_592), .ZN(n_0_0_226));
   OAI21_X1 i_0_0_478 (.A(n_0_0_227), .B1(n_0_0_236), .B2(n_0_0_474), .ZN(
      n_0_625));
   AOI222_X1 i_0_0_479 (.A1(n_0_0_241), .A2(n_0_593), .B1(n_0_86), .B2(n_0_0_238), 
      .C1(n_0_0_243), .C2(n_0_609), .ZN(n_0_0_227));
   OAI21_X1 i_0_0_480 (.A(n_0_0_228), .B1(n_0_0_236), .B2(n_0_0_475), .ZN(
      n_0_626));
   AOI222_X1 i_0_0_481 (.A1(n_0_610), .A2(n_0_0_243), .B1(n_0_0_241), .B2(
      n_0_594), .C1(n_0_87), .C2(n_0_0_238), .ZN(n_0_0_228));
   NAND2_X1 i_0_0_482 (.A1(n_0_0_229), .A2(n_0_0_230), .ZN(n_0_627));
   AOI222_X1 i_0_0_483 (.A1(n_0_88), .A2(n_0_0_238), .B1(n_0_0_237), .B2(n_0_66), 
      .C1(n_0_0_243), .C2(n_0_611), .ZN(n_0_0_229));
   NAND2_X1 i_0_0_484 (.A1(n_0_0_241), .A2(n_0_595), .ZN(n_0_0_230));
   OAI21_X1 i_0_0_485 (.A(n_0_0_231), .B1(n_0_0_236), .B2(n_0_0_66), .ZN(n_0_628));
   AOI222_X1 i_0_0_486 (.A1(n_0_0_241), .A2(n_0_596), .B1(n_0_89), .B2(n_0_0_238), 
      .C1(n_0_0_243), .C2(n_0_612), .ZN(n_0_0_231));
   OAI21_X1 i_0_0_487 (.A(n_0_0_232), .B1(n_0_0_236), .B2(n_0_0_67), .ZN(n_0_629));
   AOI222_X1 i_0_0_488 (.A1(n_0_0_241), .A2(n_0_597), .B1(n_0_90), .B2(n_0_0_238), 
      .C1(n_0_0_243), .C2(n_0_613), .ZN(n_0_0_232));
   OAI21_X1 i_0_0_489 (.A(n_0_0_233), .B1(n_0_0_236), .B2(n_0_0_68), .ZN(n_0_630));
   AOI222_X1 i_0_0_490 (.A1(n_0_614), .A2(n_0_0_243), .B1(n_0_0_241), .B2(
      n_0_598), .C1(n_0_91), .C2(n_0_0_238), .ZN(n_0_0_233));
   OAI21_X1 i_0_0_491 (.A(n_0_0_234), .B1(n_0_0_240), .B2(n_0_0_257), .ZN(
      n_0_631));
   AOI221_X1 i_0_0_492 (.A(n_0_0_239), .B1(n_0_0_238), .B2(n_0_92), .C1(
      n_0_0_237), .C2(n_0_70), .ZN(n_0_0_234));
   OAI21_X1 i_0_0_493 (.A(n_0_0_235), .B1(n_0_0_240), .B2(n_0_0_258), .ZN(
      n_0_632));
   AOI221_X1 i_0_0_494 (.A(n_0_0_239), .B1(n_0_0_238), .B2(n_0_93), .C1(
      n_0_0_237), .C2(n_0_71), .ZN(n_0_0_235));
   INV_X1 i_0_0_495 (.A(n_0_0_237), .ZN(n_0_0_236));
   NOR2_X1 i_0_0_496 (.A1(n_0_0_430), .A2(n_0_0_242), .ZN(n_0_0_237));
   NOR2_X1 i_0_0_497 (.A1(n_0_0_262), .A2(n_0_0_245), .ZN(n_0_0_238));
   NOR3_X1 i_0_0_498 (.A1(poolingReset), .A2(n_0_0_431), .A3(n_0_0_244), 
      .ZN(n_0_0_239));
   NOR2_X1 i_0_0_499 (.A1(n_0_0_243), .A2(n_0_0_241), .ZN(n_0_0_240));
   AND2_X1 i_0_0_500 (.A1(n_0_0_242), .A2(n_0_0_431), .ZN(n_0_0_241));
   NAND3_X1 i_0_0_501 (.A1(convResetState[1]), .A2(n_0_0_349), .A3(n_0_0_267), 
      .ZN(n_0_0_242));
   NOR2_X1 i_0_0_502 (.A1(n_0_0_431), .A2(n_0_0_244), .ZN(n_0_0_243));
   NOR2_X1 i_0_0_503 (.A1(n_0_0_263), .A2(n_0_0_245), .ZN(n_0_0_244));
   NAND2_X1 i_0_0_504 (.A1(poolingState[0]), .A2(n_0_0_281), .ZN(n_0_0_245));
   NAND2_X1 i_0_0_505 (.A1(poolingReset), .A2(n_0_0_247), .ZN(n_0_601));
   NAND2_X1 i_0_0_506 (.A1(poolingReset), .A2(n_0_0_248), .ZN(n_0_602));
   AND2_X1 i_0_0_507 (.A1(poolingReset), .A2(n_0_587), .ZN(n_0_603));
   MUX2_X1 i_0_0_508 (.A(writeAdress[3]), .B(n_0_0_29), .S(n_0_0_246), .Z(
      n_0_604));
   MUX2_X1 i_0_0_509 (.A(writeAdress[4]), .B(n_0_548), .S(n_0_0_246), .Z(n_0_605));
   MUX2_X1 i_0_0_510 (.A(writeAdress[5]), .B(n_0_646), .S(n_0_0_246), .Z(n_0_606));
   MUX2_X1 i_0_0_511 (.A(writeAdress[6]), .B(n_0_645), .S(n_0_0_246), .Z(n_0_607));
   MUX2_X1 i_0_0_512 (.A(writeAdress[7]), .B(n_0_0_380), .S(n_0_0_246), .Z(
      n_0_608));
   MUX2_X1 i_0_0_513 (.A(writeAdress[8]), .B(n_0_0_451), .S(n_0_0_246), .Z(
      n_0_609));
   MUX2_X1 i_0_0_514 (.A(writeAdress[9]), .B(n_0_0_253), .S(n_0_0_246), .Z(
      n_0_610));
   MUX2_X1 i_0_0_515 (.A(writeAdress[10]), .B(n_0_0_254), .S(n_0_0_246), 
      .Z(n_0_611));
   MUX2_X1 i_0_0_516 (.A(writeAdress[11]), .B(n_0_0_56), .S(n_0_0_246), .Z(
      n_0_612));
   MUX2_X1 i_0_0_517 (.A(writeAdress[12]), .B(n_0_581), .S(n_0_0_246), .Z(
      n_0_613));
   MUX2_X1 i_0_0_518 (.A(writeAdress[13]), .B(n_0_0_29), .S(n_0_0_246), .Z(
      n_0_614));
   NAND2_X1 i_0_0_519 (.A1(writeReset), .A2(poolingReset), .ZN(n_0_0_246));
   NAND2_X1 i_0_0_520 (.A1(poolingReset), .A2(n_0_0_257), .ZN(n_0_615));
   NAND2_X1 i_0_0_521 (.A1(poolingReset), .A2(n_0_0_258), .ZN(n_0_616));
   INV_X1 i_0_0_522 (.A(n_0_0_247), .ZN(n_0_585));
   NOR2_X1 i_0_0_523 (.A1(n_0_0_69), .A2(writeAdress[0]), .ZN(n_0_0_247));
   INV_X1 i_0_0_524 (.A(n_0_0_248), .ZN(n_0_586));
   NOR2_X1 i_0_0_525 (.A1(n_0_0_69), .A2(writeAdress[1]), .ZN(n_0_0_248));
   AND2_X1 i_0_0_526 (.A1(writeAdress[2]), .A2(writeReset), .ZN(n_0_587));
   MUX2_X1 i_0_0_527 (.A(writeAdress[3]), .B(n_0_0_29), .S(n_0_0_69), .Z(n_0_588));
   OAI21_X1 i_0_0_528 (.A(n_0_0_249), .B1(n_0_0_456), .B2(writeReset), .ZN(
      n_0_589));
   NAND2_X1 i_0_0_529 (.A1(writeAdress[4]), .A2(writeReset), .ZN(n_0_0_249));
   OAI21_X1 i_0_0_530 (.A(n_0_0_250), .B1(n_0_0_463), .B2(writeReset), .ZN(
      n_0_590));
   NAND2_X1 i_0_0_531 (.A1(writeAdress[5]), .A2(writeReset), .ZN(n_0_0_250));
   MUX2_X1 i_0_0_532 (.A(writeAdress[6]), .B(n_0_645), .S(n_0_0_69), .Z(n_0_591));
   OAI21_X1 i_0_0_533 (.A(n_0_0_251), .B1(n_0_0_381), .B2(writeReset), .ZN(
      n_0_592));
   NAND2_X1 i_0_0_534 (.A1(writeAdress[7]), .A2(writeReset), .ZN(n_0_0_251));
   OAI21_X1 i_0_0_535 (.A(n_0_0_252), .B1(n_0_0_450), .B2(writeReset), .ZN(
      n_0_593));
   NAND2_X1 i_0_0_536 (.A1(writeAdress[8]), .A2(writeReset), .ZN(n_0_0_252));
   MUX2_X1 i_0_0_537 (.A(writeAdress[9]), .B(n_0_0_253), .S(n_0_0_69), .Z(
      n_0_594));
   NAND2_X1 i_0_0_538 (.A1(n_0_0_461), .A2(n_0_0_442), .ZN(n_0_0_253));
   OAI21_X1 i_0_0_539 (.A(n_0_0_256), .B1(n_0_0_255), .B2(writeReset), .ZN(
      n_0_595));
   INV_X1 i_0_0_540 (.A(n_0_0_255), .ZN(n_0_0_254));
   NAND2_X1 i_0_0_541 (.A1(n_0_0_448), .A2(layerCounter[0]), .ZN(n_0_0_255));
   NAND2_X1 i_0_0_542 (.A1(writeAdress[10]), .A2(writeReset), .ZN(n_0_0_256));
   MUX2_X1 i_0_0_543 (.A(writeAdress[11]), .B(n_0_0_56), .S(n_0_0_69), .Z(
      n_0_596));
   MUX2_X1 i_0_0_544 (.A(writeAdress[12]), .B(n_0_581), .S(n_0_0_69), .Z(n_0_597));
   MUX2_X1 i_0_0_545 (.A(writeAdress[13]), .B(n_0_0_29), .S(n_0_0_69), .Z(
      n_0_598));
   INV_X1 i_0_0_546 (.A(n_0_0_257), .ZN(n_0_599));
   NOR2_X1 i_0_0_547 (.A1(n_0_0_69), .A2(writeAdress[14]), .ZN(n_0_0_257));
   INV_X1 i_0_0_548 (.A(n_0_0_258), .ZN(n_0_600));
   NOR2_X1 i_0_0_549 (.A1(n_0_0_69), .A2(writeAdress[15]), .ZN(n_0_0_258));
   NOR2_X1 i_0_0_550 (.A1(n_0_0_434), .A2(n_0_0_433), .ZN(n_0_584));
   NOR4_X1 i_0_0_558 (.A1(n_0_0_262), .A2(n_0_0_283), .A3(DMA_start), .A4(
      n_0_0_278), .ZN(n_0_0_260));
   NOR2_X1 i_0_0_559 (.A1(n_0_0_278), .A2(DMA_start), .ZN(n_0_0_261));
   OR2_X1 i_0_0_560 (.A1(n_0_0_76), .A2(n_0_0_263), .ZN(n_0_0_262));
   OR3_X1 i_0_0_561 (.A1(n_0_0_433), .A2(n_0_0_328), .A3(n_0_0_307), .ZN(
      n_0_0_263));
   NOR3_X1 i_0_0_562 (.A1(n_0_0_430), .A2(n_0_0_268), .A3(n_0_0_266), .ZN(
      n_0_0_264));
   NOR2_X1 i_0_0_563 (.A1(n_0_0_268), .A2(n_0_0_266), .ZN(n_0_0_265));
   INV_X1 i_0_0_564 (.A(n_0_0_267), .ZN(n_0_0_266));
   AND2_X1 i_0_0_565 (.A1(n_0_0_369), .A2(n_0_0_74), .ZN(n_0_0_267));
   OAI21_X1 i_0_0_566 (.A(n_0_0_70), .B1(n_0_0_350), .B2(filterCounter[31]), 
      .ZN(n_0_0_268));
   AOI211_X1 i_0_0_567 (.A(n_0_0_277), .B(n_0_0_270), .C1(n_0_0_431), .C2(
      n_0_0_397), .ZN(n_0_567));
   NAND2_X1 i_0_0_568 (.A1(n_0_0_274), .A2(n_0_0_271), .ZN(n_0_0_269));
   NOR2_X1 i_0_0_569 (.A1(n_0_0_430), .A2(n_0_0_272), .ZN(n_0_0_270));
   NOR2_X1 i_0_0_570 (.A1(n_0_0_72), .A2(n_0_0_430), .ZN(n_0_0_271));
   NAND2_X1 i_0_0_571 (.A1(convResetState[1]), .A2(n_0_0_274), .ZN(n_0_0_272));
   NOR2_X1 i_0_0_572 (.A1(n_0_0_72), .A2(n_0_0_275), .ZN(n_0_0_273));
   INV_X1 i_0_0_573 (.A(n_0_0_275), .ZN(n_0_0_274));
   OAI21_X1 i_0_0_574 (.A(n_0_0_423), .B1(n_0_0_350), .B2(filterCounter[31]), 
      .ZN(n_0_0_275));
   NAND2_X1 i_0_0_575 (.A1(n_0_0_430), .A2(n_0_0_429), .ZN(n_0_0_276));
   NOR2_X1 i_0_0_576 (.A1(n_0_0_431), .A2(n_0_0_278), .ZN(n_0_0_277));
   OR2_X1 i_0_0_577 (.A1(poolingState[1]), .A2(poolingState[0]), .ZN(n_0_0_278));
   NOR2_X1 i_0_0_579 (.A1(n_0_0_430), .A2(convResetState[1]), .ZN(n_0_568));
   NOR2_X1 i_0_0_580 (.A1(reset), .A2(n_0_0_280), .ZN(n_0_569));
   AOI21_X1 i_0_0_581 (.A(n_0_0_347), .B1(n_0_0_302), .B2(n_0_0_281), .ZN(
      n_0_0_280));
   NOR2_X1 i_0_0_582 (.A1(poolingState[1]), .A2(n_0_0_283), .ZN(n_0_0_281));
   INV_X1 i_0_0_583 (.A(n_0_0_283), .ZN(n_0_0_282));
   AOI21_X1 i_0_0_584 (.A(poolingWindowY[31]), .B1(n_0_0_284), .B2(n_0_0_285), 
      .ZN(n_0_0_283));
   AOI211_X1 i_0_0_585 (.A(n_0_0_296), .B(n_0_0_291), .C1(poolingWindowY[4]), 
      .C2(n_0_539), .ZN(n_0_0_284));
   OAI21_X1 i_0_0_586 (.A(n_0_0_286), .B1(n_0_539), .B2(poolingWindowY[4]), 
      .ZN(n_0_0_285));
   OAI22_X1 i_0_0_587 (.A1(n_0_0_287), .A2(n_0_0_395), .B1(n_0_0_290), .B2(
      n_0_0_452), .ZN(n_0_0_286));
   AOI22_X1 i_0_0_588 (.A1(n_0_0_288), .A2(poolingWindowY[2]), .B1(
      poolingWindowY[1]), .B2(n_0_0_451), .ZN(n_0_0_287));
   NAND2_X1 i_0_0_589 (.A1(n_0_0_453), .A2(n_0_0_289), .ZN(n_0_0_288));
   NAND2_X1 i_0_0_590 (.A1(poolingWindowY[1]), .A2(n_0_0_460), .ZN(n_0_0_289));
   NOR3_X1 i_0_0_591 (.A1(n_0_0_65), .A2(poolingWindowY[2]), .A3(
      poolingWindowY[3]), .ZN(n_0_0_290));
   NAND4_X1 i_0_0_592 (.A1(n_0_0_295), .A2(n_0_0_294), .A3(n_0_0_293), .A4(
      n_0_0_292), .ZN(n_0_0_291));
   NOR4_X1 i_0_0_593 (.A1(poolingWindowY[30]), .A2(poolingWindowY[29]), .A3(
      poolingWindowY[28]), .A4(poolingWindowY[27]), .ZN(n_0_0_292));
   NOR4_X1 i_0_0_594 (.A1(poolingWindowY[26]), .A2(poolingWindowY[25]), .A3(
      poolingWindowY[24]), .A4(poolingWindowY[17]), .ZN(n_0_0_293));
   NOR2_X1 i_0_0_595 (.A1(poolingWindowY[23]), .A2(poolingWindowY[22]), .ZN(
      n_0_0_294));
   NOR4_X1 i_0_0_596 (.A1(poolingWindowY[21]), .A2(poolingWindowY[20]), .A3(
      poolingWindowY[19]), .A4(poolingWindowY[18]), .ZN(n_0_0_295));
   NAND4_X1 i_0_0_597 (.A1(n_0_0_300), .A2(n_0_0_299), .A3(n_0_0_298), .A4(
      n_0_0_297), .ZN(n_0_0_296));
   NOR4_X1 i_0_0_598 (.A1(poolingWindowY[16]), .A2(poolingWindowY[11]), .A3(
      poolingWindowY[9]), .A4(poolingWindowY[8]), .ZN(n_0_0_297));
   NOR2_X1 i_0_0_599 (.A1(poolingWindowY[10]), .A2(poolingWindowY[7]), .ZN(
      n_0_0_298));
   NOR2_X1 i_0_0_600 (.A1(poolingWindowY[6]), .A2(poolingWindowY[5]), .ZN(
      n_0_0_299));
   AND2_X1 i_0_0_601 (.A1(n_0_0_301), .A2(n_0_0_436), .ZN(n_0_0_300));
   NOR4_X1 i_0_0_602 (.A1(poolingWindowY[15]), .A2(poolingWindowY[14]), .A3(
      poolingWindowY[13]), .A4(poolingWindowY[12]), .ZN(n_0_0_301));
   INV_X1 i_0_0_603 (.A(n_0_0_303), .ZN(n_0_0_302));
   OR2_X1 i_0_0_604 (.A1(n_0_0_304), .A2(n_0_0_328), .ZN(n_0_0_303));
   NAND3_X1 i_0_0_605 (.A1(n_0_0_306), .A2(n_0_0_427), .A3(layerCounter[0]), 
      .ZN(n_0_0_304));
   NAND2_X1 i_0_0_606 (.A1(layerCounter[0]), .A2(n_0_0_427), .ZN(n_0_0_305));
   INV_X1 i_0_0_607 (.A(n_0_0_307), .ZN(n_0_0_306));
   NOR2_X1 i_0_0_608 (.A1(poolingCounter[31]), .A2(n_0_0_308), .ZN(n_0_0_307));
   NOR4_X1 i_0_0_609 (.A1(n_0_0_309), .A2(n_0_0_318), .A3(n_0_0_323), .A4(
      n_0_0_316), .ZN(n_0_0_308));
   AOI22_X1 i_0_0_610 (.A1(n_0_0_314), .A2(n_0_0_312), .B1(n_0_0_310), .B2(
      n_0_0_61), .ZN(n_0_0_309));
   OAI21_X1 i_0_0_611 (.A(poolingCounter[4]), .B1(n_0_0_445), .B2(n_0_0_311), 
      .ZN(n_0_0_310));
   AND2_X1 i_0_0_612 (.A1(poolingCounter[6]), .A2(poolingCounter[5]), .ZN(
      n_0_0_311));
   OAI21_X1 i_0_0_613 (.A(n_0_0_76), .B1(n_0_0_313), .B2(layerCounter[2]), 
      .ZN(n_0_0_312));
   AOI21_X1 i_0_0_614 (.A(layerCounter[1]), .B1(n_0_0_259), .B2(n_0_0_279), 
      .ZN(n_0_0_313));
   AOI221_X1 i_0_0_615 (.A(poolingCounter[3]), .B1(layerCounter[1]), .B2(
      layerCounter[0]), .C1(n_0_0_315), .C2(poolingCounter[2]), .ZN(n_0_0_314));
   OAI21_X1 i_0_0_616 (.A(n_0_0_65), .B1(layerCounter[2]), .B2(n_0_0_279), 
      .ZN(n_0_0_315));
   INV_X1 i_0_0_617 (.A(n_0_0_317), .ZN(n_0_0_316));
   OAI21_X1 i_0_0_618 (.A(n_0_0_445), .B1(poolingCounter[5]), .B2(
      poolingCounter[6]), .ZN(n_0_0_317));
   NAND4_X1 i_0_0_619 (.A1(n_0_0_322), .A2(n_0_0_321), .A3(n_0_0_320), .A4(
      n_0_0_319), .ZN(n_0_0_318));
   NOR4_X1 i_0_0_620 (.A1(poolingCounter[31]), .A2(poolingCounter[30]), .A3(
      poolingCounter[29]), .A4(poolingCounter[28]), .ZN(n_0_0_319));
   NOR4_X1 i_0_0_621 (.A1(poolingCounter[27]), .A2(poolingCounter[26]), .A3(
      poolingCounter[25]), .A4(poolingCounter[18]), .ZN(n_0_0_320));
   NOR4_X1 i_0_0_622 (.A1(poolingCounter[23]), .A2(poolingCounter[22]), .A3(
      poolingCounter[21]), .A4(poolingCounter[20]), .ZN(n_0_0_321));
   NOR2_X1 i_0_0_623 (.A1(poolingCounter[24]), .A2(poolingCounter[19]), .ZN(
      n_0_0_322));
   NAND4_X1 i_0_0_624 (.A1(n_0_0_327), .A2(n_0_0_326), .A3(n_0_0_325), .A4(
      n_0_0_324), .ZN(n_0_0_323));
   NOR3_X1 i_0_0_625 (.A1(poolingCounter[16]), .A2(poolingCounter[15]), .A3(
      poolingCounter[14]), .ZN(n_0_0_324));
   NOR4_X1 i_0_0_626 (.A1(poolingCounter[17]), .A2(poolingCounter[13]), .A3(
      poolingCounter[12]), .A4(poolingCounter[10]), .ZN(n_0_0_325));
   NOR4_X1 i_0_0_627 (.A1(poolingCounter[11]), .A2(poolingCounter[9]), .A3(
      poolingCounter[8]), .A4(poolingCounter[7]), .ZN(n_0_0_326));
   NAND3_X1 i_0_0_628 (.A1(n_0_0_450), .A2(n_0_0_448), .A3(poolingCounter[4]), 
      .ZN(n_0_0_327));
   AOI21_X1 i_0_0_629 (.A(poolingWindowX[31]), .B1(n_0_0_329), .B2(n_0_0_330), 
      .ZN(n_0_0_328));
   AOI211_X1 i_0_0_630 (.A(n_0_0_341), .B(n_0_0_336), .C1(poolingWindowX[4]), 
      .C2(n_0_539), .ZN(n_0_0_329));
   OAI21_X1 i_0_0_631 (.A(n_0_0_331), .B1(n_0_539), .B2(poolingWindowX[4]), 
      .ZN(n_0_0_330));
   OAI22_X1 i_0_0_632 (.A1(n_0_0_332), .A2(n_0_0_393), .B1(n_0_0_335), .B2(
      n_0_0_452), .ZN(n_0_0_331));
   AOI22_X1 i_0_0_633 (.A1(n_0_0_333), .A2(poolingWindowX[2]), .B1(
      poolingWindowX[1]), .B2(n_0_0_451), .ZN(n_0_0_332));
   NAND2_X1 i_0_0_634 (.A1(n_0_0_453), .A2(n_0_0_334), .ZN(n_0_0_333));
   NAND2_X1 i_0_0_635 (.A1(poolingWindowX[1]), .A2(n_0_0_460), .ZN(n_0_0_334));
   NOR3_X1 i_0_0_636 (.A1(n_0_0_65), .A2(poolingWindowX[2]), .A3(
      poolingWindowX[3]), .ZN(n_0_0_335));
   NAND4_X1 i_0_0_637 (.A1(n_0_0_340), .A2(n_0_0_339), .A3(n_0_0_338), .A4(
      n_0_0_337), .ZN(n_0_0_336));
   NOR4_X1 i_0_0_638 (.A1(poolingWindowX[30]), .A2(poolingWindowX[29]), .A3(
      poolingWindowX[28]), .A4(poolingWindowX[27]), .ZN(n_0_0_337));
   NOR4_X1 i_0_0_639 (.A1(poolingWindowX[26]), .A2(poolingWindowX[25]), .A3(
      poolingWindowX[24]), .A4(poolingWindowX[17]), .ZN(n_0_0_338));
   NOR2_X1 i_0_0_640 (.A1(poolingWindowX[23]), .A2(poolingWindowX[22]), .ZN(
      n_0_0_339));
   NOR4_X1 i_0_0_641 (.A1(poolingWindowX[21]), .A2(poolingWindowX[20]), .A3(
      poolingWindowX[19]), .A4(poolingWindowX[18]), .ZN(n_0_0_340));
   NAND4_X1 i_0_0_642 (.A1(n_0_0_345), .A2(n_0_0_344), .A3(n_0_0_343), .A4(
      n_0_0_342), .ZN(n_0_0_341));
   NOR4_X1 i_0_0_643 (.A1(poolingWindowX[16]), .A2(poolingWindowX[11]), .A3(
      poolingWindowX[9]), .A4(poolingWindowX[8]), .ZN(n_0_0_342));
   NOR2_X1 i_0_0_644 (.A1(poolingWindowX[10]), .A2(poolingWindowX[7]), .ZN(
      n_0_0_343));
   NOR2_X1 i_0_0_645 (.A1(poolingWindowX[6]), .A2(poolingWindowX[5]), .ZN(
      n_0_0_344));
   AND2_X1 i_0_0_646 (.A1(n_0_0_346), .A2(n_0_0_436), .ZN(n_0_0_345));
   NOR4_X1 i_0_0_647 (.A1(poolingWindowX[15]), .A2(poolingWindowX[14]), .A3(
      poolingWindowX[13]), .A4(poolingWindowX[12]), .ZN(n_0_0_346));
   AOI211_X1 i_0_0_648 (.A(layerCounter[0]), .B(n_0_0_426), .C1(n_0_0_348), 
      .C2(convResetState[1]), .ZN(n_0_0_347));
   OAI21_X1 i_0_0_649 (.A(n_0_0_369), .B1(n_0_0_349), .B2(n_0_0_70), .ZN(
      n_0_0_348));
   NOR2_X1 i_0_0_650 (.A1(filterCounter[31]), .A2(n_0_0_350), .ZN(n_0_0_349));
   INV_X1 i_0_0_651 (.A(n_0_0_351), .ZN(n_0_0_350));
   OAI21_X1 i_0_0_652 (.A(n_0_0_357), .B1(n_0_0_352), .B2(n_0_0_446), .ZN(
      n_0_0_351));
   NOR4_X1 i_0_0_653 (.A1(filterCounter[6]), .A2(filterCounter[5]), .A3(
      filterCounter[4]), .A4(n_0_0_353), .ZN(n_0_0_352));
   NOR3_X1 i_0_0_654 (.A1(n_0_0_354), .A2(n_0_0_28), .A3(n_0_0_355), .ZN(
      n_0_0_353));
   AOI211_X1 i_0_0_655 (.A(filterCounter[3]), .B(n_0_0_463), .C1(
      filterCounter[1]), .C2(filterCounter[2]), .ZN(n_0_0_354));
   NOR4_X1 i_0_0_656 (.A1(n_0_0_356), .A2(filterCounter[0]), .A3(
      filterCounter[1]), .A4(filterCounter[2]), .ZN(n_0_0_355));
   OR2_X1 i_0_0_657 (.A1(n_0_0_65), .A2(filterCounter[3]), .ZN(n_0_0_356));
   NOR3_X1 i_0_0_658 (.A1(n_0_0_364), .A2(n_0_0_361), .A3(n_0_0_358), .ZN(
      n_0_0_357));
   NAND2_X1 i_0_0_659 (.A1(n_0_0_360), .A2(n_0_0_359), .ZN(n_0_0_358));
   NOR4_X1 i_0_0_660 (.A1(filterCounter[28]), .A2(filterCounter[27]), .A3(
      filterCounter[26]), .A4(filterCounter[25]), .ZN(n_0_0_359));
   NOR4_X1 i_0_0_661 (.A1(filterCounter[30]), .A2(filterCounter[29]), .A3(
      filterCounter[10]), .A4(filterCounter[7]), .ZN(n_0_0_360));
   NAND3_X1 i_0_0_662 (.A1(n_0_0_368), .A2(n_0_0_363), .A3(n_0_0_362), .ZN(
      n_0_0_361));
   NOR2_X1 i_0_0_663 (.A1(filterCounter[23]), .A2(filterCounter[18]), .ZN(
      n_0_0_362));
   NOR4_X1 i_0_0_664 (.A1(filterCounter[24]), .A2(filterCounter[22]), .A3(
      filterCounter[21]), .A4(filterCounter[17]), .ZN(n_0_0_363));
   NAND3_X1 i_0_0_665 (.A1(n_0_0_366), .A2(n_0_0_365), .A3(n_0_0_367), .ZN(
      n_0_0_364));
   NOR4_X1 i_0_0_666 (.A1(filterCounter[16]), .A2(filterCounter[11]), .A3(
      filterCounter[9]), .A4(filterCounter[8]), .ZN(n_0_0_365));
   NOR4_X1 i_0_0_667 (.A1(filterCounter[15]), .A2(filterCounter[14]), .A3(
      filterCounter[13]), .A4(filterCounter[12]), .ZN(n_0_0_366));
   NAND4_X1 i_0_0_668 (.A1(filterCounter[6]), .A2(filterCounter[5]), .A3(
      filterCounter[4]), .A4(filterCounter[3]), .ZN(n_0_0_367));
   NOR2_X1 i_0_0_669 (.A1(filterCounter[20]), .A2(filterCounter[19]), .ZN(
      n_0_0_368));
   NOR3_X1 i_0_0_670 (.A1(n_0_0_424), .A2(n_0_0_389), .A3(n_0_0_372), .ZN(
      n_0_0_369));
   NOR2_X1 i_0_0_671 (.A1(n_0_0_424), .A2(n_0_0_389), .ZN(n_0_0_370));
   INV_X1 i_0_0_672 (.A(n_0_0_372), .ZN(n_0_0_371));
   AOI21_X1 i_0_0_673 (.A(kernelCounter[31]), .B1(n_0_0_382), .B2(n_0_0_373), 
      .ZN(n_0_0_372));
   AOI21_X1 i_0_0_674 (.A(n_0_0_374), .B1(n_0_0_378), .B2(kernelCounter[3]), 
      .ZN(n_0_0_373));
   NAND4_X1 i_0_0_675 (.A1(n_0_0_57), .A2(n_0_0_377), .A3(n_0_0_376), .A4(
      n_0_0_375), .ZN(n_0_0_374));
   NAND4_X1 i_0_0_676 (.A1(n_0_0_86), .A2(n_0_0_85), .A3(kernelCounter[2]), 
      .A4(kernelCounter[1]), .ZN(n_0_0_375));
   NOR4_X1 i_0_0_677 (.A1(kernelCounter[13]), .A2(kernelCounter[12]), .A3(
      kernelCounter[11]), .A4(kernelCounter[10]), .ZN(n_0_0_376));
   NOR4_X1 i_0_0_679 (.A1(kernelCounter[28]), .A2(kernelCounter[14]), .A3(
      kernelCounter[9]), .A4(kernelCounter[7]), .ZN(n_0_0_377));
   NAND2_X1 i_0_0_680 (.A1(n_0_0_380), .A2(n_0_0_379), .ZN(n_0_0_378));
   NAND3_X1 i_0_0_681 (.A1(kernelCounter[6]), .A2(kernelCounter[5]), .A3(
      kernelCounter[4]), .ZN(n_0_0_379));
   INV_X1 i_0_0_682 (.A(n_0_0_381), .ZN(n_0_0_380));
   NAND2_X1 i_0_0_683 (.A1(n_0_0_57), .A2(n_0_0_454), .ZN(n_0_0_381));
   AOI21_X1 i_0_0_684 (.A(n_0_0_384), .B1(n_0_0_383), .B2(n_0_0_462), .ZN(
      n_0_0_382));
   OR3_X1 i_0_0_685 (.A1(kernelCounter[6]), .A2(kernelCounter[5]), .A3(
      kernelCounter[4]), .ZN(n_0_0_383));
   NAND4_X1 i_0_0_686 (.A1(n_0_0_388), .A2(n_0_0_387), .A3(n_0_0_386), .A4(
      n_0_0_385), .ZN(n_0_0_384));
   NOR4_X1 i_0_0_687 (.A1(kernelCounter[22]), .A2(kernelCounter[20]), .A3(
      kernelCounter[19]), .A4(kernelCounter[15]), .ZN(n_0_0_385));
   NOR4_X1 i_0_0_688 (.A1(kernelCounter[21]), .A2(kernelCounter[18]), .A3(
      kernelCounter[17]), .A4(kernelCounter[16]), .ZN(n_0_0_386));
   NOR4_X1 i_0_0_689 (.A1(kernelCounter[30]), .A2(kernelCounter[29]), .A3(
      kernelCounter[27]), .A4(kernelCounter[8]), .ZN(n_0_0_387));
   NOR4_X1 i_0_0_690 (.A1(kernelCounter[26]), .A2(kernelCounter[25]), .A3(
      kernelCounter[24]), .A4(kernelCounter[23]), .ZN(n_0_0_388));
   AOI22_X1 i_0_0_691 (.A1(n_0_0_407), .A2(n_0_0_404), .B1(n_0_0_390), .B2(
      convWindowX[31]), .ZN(n_0_0_389));
   NAND2_X1 i_0_0_692 (.A1(n_0_0_400), .A2(n_0_0_391), .ZN(n_0_0_390));
   NOR4_X1 i_0_0_693 (.A1(n_0_0_399), .A2(n_0_0_398), .A3(n_0_0_394), .A4(
      n_0_0_392), .ZN(n_0_0_391));
   NAND4_X1 i_0_0_694 (.A1(convWindowX[30]), .A2(convWindowX[29]), .A3(
      convWindowX[28]), .A4(convWindowX[27]), .ZN(n_0_0_392));
   NAND4_X1 i_0_0_695 (.A1(convWindowX[26]), .A2(convWindowX[25]), .A3(
      convWindowX[24]), .A4(convWindowX[17]), .ZN(n_0_0_394));
   NAND4_X1 i_0_0_696 (.A1(convWindowX[22]), .A2(convWindowX[21]), .A3(
      convWindowX[20]), .A4(convWindowX[19]), .ZN(n_0_0_398));
   NAND2_X1 i_0_0_697 (.A1(convWindowX[23]), .A2(convWindowX[18]), .ZN(n_0_0_399));
   NOR4_X1 i_0_0_698 (.A1(n_0_0_423), .A2(n_0_0_403), .A3(n_0_0_402), .A4(
      n_0_0_401), .ZN(n_0_0_400));
   NAND4_X1 i_0_0_699 (.A1(convWindowX[16]), .A2(convWindowX[11]), .A3(
      convWindowX[9]), .A4(convWindowX[8]), .ZN(n_0_0_401));
   NAND4_X1 i_0_0_700 (.A1(convWindowX[10]), .A2(convWindowX[7]), .A3(
      convWindowX[6]), .A4(convWindowX[5]), .ZN(n_0_0_402));
   NAND4_X1 i_0_0_701 (.A1(convWindowX[15]), .A2(convWindowX[14]), .A3(
      convWindowX[13]), .A4(convWindowX[12]), .ZN(n_0_0_403));
   OAI21_X1 i_0_0_702 (.A(convWindowX[3]), .B1(n_0_0_405), .B2(n_0_0_28), 
      .ZN(n_0_0_404));
   AOI21_X1 i_0_0_703 (.A(n_0_0_396), .B1(n_0_0_453), .B2(n_0_0_406), .ZN(
      n_0_0_405));
   OAI21_X1 i_0_0_704 (.A(convWindowX[2]), .B1(n_0_0_410), .B2(n_0_0_458), 
      .ZN(n_0_0_406));
   AOI221_X1 i_0_0_705 (.A(n_0_0_413), .B1(n_0_0_410), .B2(n_0_0_408), .C1(
      n_0_0_29), .C2(convWindowX[4]), .ZN(n_0_0_407));
   OAI21_X1 i_0_0_706 (.A(n_0_0_462), .B1(n_0_0_456), .B2(n_0_0_409), .ZN(
      n_0_0_408));
   AOI21_X1 i_0_0_707 (.A(convWindowX[3]), .B1(convWindowX[2]), .B2(
      layerCounter[0]), .ZN(n_0_0_409));
   NAND2_X1 i_0_0_708 (.A1(n_0_0_412), .A2(n_0_0_411), .ZN(n_0_0_410));
   AOI21_X1 i_0_0_709 (.A(convWindowX[1]), .B1(convWindowX[0]), .B2(
      layerCounter[2]), .ZN(n_0_0_411));
   NAND2_X1 i_0_0_710 (.A1(convWindowX[2]), .A2(n_0_0_57), .ZN(n_0_0_412));
   AOI21_X1 i_0_0_711 (.A(convWindowX[31]), .B1(n_0_0_419), .B2(n_0_0_414), 
      .ZN(n_0_0_413));
   AND4_X1 i_0_0_712 (.A1(n_0_0_418), .A2(n_0_0_417), .A3(n_0_0_416), .A4(
      n_0_0_415), .ZN(n_0_0_414));
   NOR4_X1 i_0_0_713 (.A1(convWindowX[30]), .A2(convWindowX[29]), .A3(
      convWindowX[28]), .A4(convWindowX[27]), .ZN(n_0_0_415));
   NOR4_X1 i_0_0_714 (.A1(convWindowX[26]), .A2(convWindowX[25]), .A3(
      convWindowX[24]), .A4(convWindowX[17]), .ZN(n_0_0_416));
   NOR4_X1 i_0_0_715 (.A1(convWindowX[22]), .A2(convWindowX[21]), .A3(
      convWindowX[20]), .A4(convWindowX[19]), .ZN(n_0_0_417));
   NOR2_X1 i_0_0_716 (.A1(convWindowX[23]), .A2(convWindowX[18]), .ZN(n_0_0_418));
   AND4_X1 i_0_0_717 (.A1(n_0_0_422), .A2(n_0_0_421), .A3(n_0_0_420), .A4(
      n_0_0_423), .ZN(n_0_0_419));
   NOR4_X1 i_0_0_718 (.A1(convWindowX[16]), .A2(convWindowX[11]), .A3(
      convWindowX[9]), .A4(convWindowX[8]), .ZN(n_0_0_420));
   NOR4_X1 i_0_0_719 (.A1(convWindowX[10]), .A2(convWindowX[7]), .A3(
      convWindowX[6]), .A4(convWindowX[5]), .ZN(n_0_0_421));
   NOR4_X1 i_0_0_720 (.A1(convWindowX[15]), .A2(convWindowX[14]), .A3(
      convWindowX[13]), .A4(convWindowX[12]), .ZN(n_0_0_422));
   NAND2_X1 i_0_0_721 (.A1(n_0_0_65), .A2(layerCounter[2]), .ZN(n_0_0_423));
   NOR2_X1 i_0_0_722 (.A1(n_0_0_464), .A2(n_0_0_86), .ZN(n_0_0_424));
   NOR2_X1 i_0_0_736 (.A1(n_0_0_426), .A2(layerCounter[0]), .ZN(n_0_0_425));
   NAND3_X1 i_0_0_737 (.A1(n_0_0_74), .A2(n_0_0_432), .A3(start), .ZN(n_0_0_426));
   NOR2_X1 i_0_0_738 (.A1(n_0_0_433), .A2(n_0_0_435), .ZN(n_0_0_427));
   NOR3_X1 i_0_0_739 (.A1(n_0_0_434), .A2(n_0_0_430), .A3(n_0_0_428), .ZN(
      n_0_573));
   OR2_X1 i_0_0_740 (.A1(convResetState[1]), .A2(convResetState[0]), .ZN(
      n_0_0_428));
   NAND2_X1 i_0_0_742 (.A1(n_0_0_76), .A2(n_0_0_432), .ZN(n_0_0_430));
   NOR2_X1 i_0_0_743 (.A1(layerCounter[0]), .A2(n_0_0_433), .ZN(n_0_0_431));
   INV_X1 i_0_0_744 (.A(n_0_0_433), .ZN(n_0_0_432));
   NOR2_X1 i_0_0_745 (.A1(n_0_0_465), .A2(layerCounter[31]), .ZN(n_0_0_433));
   INV_X1 i_0_0_746 (.A(n_0_0_434), .ZN(n_0_549));
   NAND3_X1 i_0_0_747 (.A1(n_0_0_74), .A2(n_0_0_73), .A3(start), .ZN(n_0_0_434));
   NAND2_X1 i_0_0_748 (.A1(n_0_0_74), .A2(start), .ZN(n_0_0_435));
   AOI21_X1 i_0_0_749 (.A(n_0_572), .B1(n_0_0_456), .B2(n_0_0_452), .ZN(n_0_540));
   NAND2_X1 i_0_0_750 (.A1(n_0_0_456), .A2(n_0_0_452), .ZN(n_0_539));
   AND2_X1 i_0_0_751 (.A1(n_0_0_65), .A2(n_0_0_436), .ZN(n_0_541));
   NAND3_X1 i_0_0_752 (.A1(layerCounter[2]), .A2(layerCounter[1]), .A3(
      layerCounter[0]), .ZN(n_0_0_436));
   AND2_X1 i_0_0_753 (.A1(n_0_0_441), .A2(n_0_0_437), .ZN(n_0_542));
   OAI21_X1 i_0_0_754 (.A(n_0_639), .B1(n_0_646), .B2(n_0_644), .ZN(n_0_0_437));
   XOR2_X1 i_0_0_755 (.A(n_0_640), .B(n_0_0_441), .Z(n_0_543));
   XNOR2_X1 i_0_0_756 (.A(n_0_641), .B(n_0_0_440), .ZN(n_0_544));
   XNOR2_X1 i_0_0_757 (.A(n_0_642), .B(n_0_0_439), .ZN(n_0_545));
   NOR2_X1 i_0_0_758 (.A1(n_0_581), .A2(n_0_0_438), .ZN(n_0_546));
   INV_X1 i_0_0_759 (.A(n_0_0_27), .ZN(n_0_547));
   XNOR2_X1 i_0_0_760 (.A(n_0_0_442), .B(n_0_0_438), .ZN(n_0_0_27));
   NOR4_X1 i_0_0_761 (.A1(n_0_0_441), .A2(n_0_640), .A3(n_0_641), .A4(n_0_642), 
      .ZN(n_0_0_438));
   NOR3_X1 i_0_0_762 (.A1(n_0_0_441), .A2(n_0_640), .A3(n_0_641), .ZN(n_0_0_439));
   NOR2_X1 i_0_0_763 (.A1(n_0_0_441), .A2(n_0_640), .ZN(n_0_0_440));
   OR3_X1 i_0_0_764 (.A1(n_0_639), .A2(n_0_646), .A3(n_0_644), .ZN(n_0_0_441));
   INV_X1 i_0_0_765 (.A(n_0_0_442), .ZN(n_0_570));
   NAND2_X1 i_0_0_766 (.A1(n_0_0_464), .A2(n_0_0_86), .ZN(n_0_0_442));
   AND2_X1 i_0_0_767 (.A1(poolingReset), .A2(readAdress[0]), .ZN(n_0_681));
   NAND2_X1 i_0_0_768 (.A1(n_0_0_466), .A2(poolingReset), .ZN(n_0_682));
   AND2_X1 i_0_0_769 (.A1(poolingReset), .A2(readAdress[2]), .ZN(n_0_683));
   MUX2_X1 i_0_0_770 (.A(n_0_0_61), .B(readAdress[3]), .S(poolingReset), 
      .Z(n_0_684));
   MUX2_X1 i_0_0_771 (.A(n_0_0_28), .B(readAdress[4]), .S(poolingReset), 
      .Z(n_0_685));
   NAND2_X1 i_0_0_772 (.A1(n_0_0_462), .A2(n_0_0_450), .ZN(n_0_0_28));
   MUX2_X1 i_0_0_773 (.A(n_0_0_29), .B(readAdress[5]), .S(poolingReset), 
      .Z(n_0_686));
   NAND2_X1 i_0_0_774 (.A1(n_0_0_462), .A2(n_0_0_456), .ZN(n_0_0_29));
   MUX2_X1 i_0_0_775 (.A(n_0_0_30), .B(readAdress[6]), .S(poolingReset), 
      .Z(n_0_687));
   NAND2_X1 i_0_0_776 (.A1(n_0_0_456), .A2(n_0_0_445), .ZN(n_0_0_30));
   MUX2_X1 i_0_0_777 (.A(n_0_0_55), .B(readAdress[7]), .S(poolingReset), 
      .Z(n_0_688));
   NAND2_X1 i_0_0_778 (.A1(n_0_0_450), .A2(n_0_0_445), .ZN(n_0_0_55));
   OAI21_X1 i_0_0_779 (.A(n_0_0_443), .B1(n_0_0_462), .B2(poolingReset), 
      .ZN(n_0_689));
   NAND2_X1 i_0_0_780 (.A1(poolingReset), .A2(readAdress[8]), .ZN(n_0_0_443));
   MUX2_X1 i_0_0_781 (.A(n_0_0_56), .B(readAdress[9]), .S(poolingReset), 
      .Z(n_0_690));
   AOI21_X1 i_0_0_782 (.A(layerCounter[1]), .B1(layerCounter[0]), .B2(
      layerCounter[2]), .ZN(n_0_0_56));
   MUX2_X1 i_0_0_783 (.A(n_0_0_57), .B(readAdress[10]), .S(poolingReset), 
      .Z(n_0_691));
   AOI21_X1 i_0_0_784 (.A(layerCounter[0]), .B1(layerCounter[1]), .B2(
      layerCounter[2]), .ZN(n_0_0_57));
   MUX2_X1 i_0_0_785 (.A(n_0_0_444), .B(readAdress[11]), .S(poolingReset), 
      .Z(n_0_692));
   INV_X1 i_0_0_786 (.A(n_0_0_444), .ZN(n_0_0_58));
   NAND2_X1 i_0_0_787 (.A1(n_0_0_457), .A2(n_0_0_445), .ZN(n_0_0_444));
   NAND2_X1 i_0_0_788 (.A1(layerCounter[0]), .A2(n_0_0_449), .ZN(n_0_0_445));
   NOR2_X1 i_0_0_789 (.A1(n_0_0_76), .A2(n_0_0_448), .ZN(n_0_0_446));
   OAI21_X1 i_0_0_790 (.A(n_0_0_447), .B1(n_0_0_455), .B2(poolingReset), 
      .ZN(n_0_693));
   NAND2_X1 i_0_0_791 (.A1(poolingReset), .A2(readAdress[12]), .ZN(n_0_0_447));
   MUX2_X1 i_0_0_792 (.A(n_0_0_61), .B(readAdress[13]), .S(poolingReset), 
      .Z(n_0_694));
   NAND2_X1 i_0_0_793 (.A1(n_0_0_450), .A2(n_0_0_448), .ZN(n_0_0_61));
   NAND2_X1 i_0_0_794 (.A1(n_0_0_85), .A2(layerCounter[2]), .ZN(n_0_0_448));
   NOR2_X1 i_0_0_795 (.A1(n_0_0_86), .A2(layerCounter[1]), .ZN(n_0_0_449));
   NAND2_X1 i_0_0_796 (.A1(layerCounter[0]), .A2(n_0_548), .ZN(n_0_0_450));
   NOR2_X1 i_0_0_797 (.A1(n_0_0_461), .A2(layerCounter[2]), .ZN(n_0_0_451));
   NAND2_X1 i_0_0_801 (.A1(n_0_0_467), .A2(poolingReset), .ZN(n_0_695));
   NAND2_X1 i_0_0_802 (.A1(n_0_0_468), .A2(poolingReset), .ZN(n_0_696));
   INV_X1 i_0_0_803 (.A(n_0_0_452), .ZN(n_0_644));
   NAND2_X1 i_0_0_804 (.A1(n_0_0_461), .A2(layerCounter[2]), .ZN(n_0_0_452));
   NAND2_X1 i_0_0_805 (.A1(n_0_0_462), .A2(n_0_0_457), .ZN(n_0_645));
   OAI21_X1 i_0_0_806 (.A(n_0_0_462), .B1(n_0_0_453), .B2(layerCounter[1]), 
      .ZN(n_0_583));
   NOR2_X1 i_0_0_807 (.A1(n_0_0_453), .A2(layerCounter[1]), .ZN(n_0_581));
   NAND2_X1 i_0_0_808 (.A1(n_0_0_86), .A2(layerCounter[0]), .ZN(n_0_0_453));
   NAND2_X1 i_0_0_809 (.A1(n_0_0_86), .A2(n_0_0_85), .ZN(n_0_0_454));
   INV_X1 i_0_0_810 (.A(n_0_0_455), .ZN(n_0_571));
   NAND2_X1 i_0_0_811 (.A1(n_0_548), .A2(n_0_0_76), .ZN(n_0_0_455));
   INV_X1 i_0_0_812 (.A(n_0_0_456), .ZN(n_0_548));
   NAND2_X1 i_0_0_813 (.A1(n_0_0_86), .A2(layerCounter[1]), .ZN(n_0_0_456));
   INV_X1 i_0_0_814 (.A(n_0_0_457), .ZN(n_0_0_62));
   NAND2_X1 i_0_0_815 (.A1(n_0_646), .A2(n_0_0_461), .ZN(n_0_0_457));
   NOR2_X1 i_0_0_816 (.A1(n_0_0_460), .A2(n_0_0_459), .ZN(n_0_0_458));
   NOR2_X1 i_0_0_817 (.A1(n_0_0_76), .A2(layerCounter[1]), .ZN(n_0_0_459));
   NOR2_X1 i_0_0_818 (.A1(n_0_0_85), .A2(layerCounter[0]), .ZN(n_0_0_460));
   NAND2_X1 i_0_0_819 (.A1(layerCounter[1]), .A2(layerCounter[0]), .ZN(n_0_0_461));
   INV_X1 i_0_0_820 (.A(n_0_0_462), .ZN(n_0_572));
   NAND2_X1 i_0_0_821 (.A1(layerCounter[2]), .A2(n_0_0_464), .ZN(n_0_0_462));
   INV_X1 i_0_0_822 (.A(n_0_0_463), .ZN(n_0_646));
   NAND2_X1 i_0_0_823 (.A1(n_0_0_86), .A2(n_0_0_65), .ZN(n_0_0_463));
   INV_X1 i_0_0_824 (.A(n_0_0_464), .ZN(n_0_0_65));
   NOR2_X1 i_0_0_825 (.A1(layerCounter[1]), .A2(layerCounter[0]), .ZN(n_0_0_464));
   INV_X1 i_0_0_826 (.A(n_0_0_1), .ZN(n_0_0_465));
   INV_X1 i_0_0_827 (.A(readAdress[1]), .ZN(n_0_0_466));
   INV_X1 i_0_0_828 (.A(readAdress[14]), .ZN(n_0_0_467));
   INV_X1 i_0_0_829 (.A(readAdress[15]), .ZN(n_0_0_468));
   INV_X1 i_0_0_830 (.A(convReset), .ZN(n_0_0_469));
   INV_X1 i_0_0_831 (.A(n_0_59), .ZN(n_0_0_470));
   INV_X1 i_0_0_832 (.A(n_0_60), .ZN(n_0_0_471));
   INV_X1 i_0_0_833 (.A(n_0_61), .ZN(n_0_0_472));
   INV_X1 i_0_0_834 (.A(n_0_62), .ZN(n_0_0_473));
   INV_X1 i_0_0_835 (.A(n_0_64), .ZN(n_0_0_474));
   INV_X1 i_0_0_836 (.A(n_0_65), .ZN(n_0_0_475));
   INV_X1 i_0_0_837 (.A(n_0_67), .ZN(n_0_0_66));
   INV_X1 i_0_0_838 (.A(n_0_68), .ZN(n_0_0_67));
   INV_X1 i_0_0_839 (.A(n_0_69), .ZN(n_0_0_68));
   INV_X1 i_0_0_840 (.A(writeReset), .ZN(n_0_0_69));
   INV_X1 i_0_0_841 (.A(convState), .ZN(n_0_0_70));
   INV_X1 i_0_0_842 (.A(poolingState[1]), .ZN(n_0_0_71));
   INV_X1 i_0_0_843 (.A(convResetState[1]), .ZN(n_0_0_72));
   INV_X1 i_0_0_844 (.A(reset), .ZN(n_0_0_73));
   INV_X1 i_0_0_856 (.A(DMA_start), .ZN(n_0_0_74));
   INV_X1 i_0_0_857 (.A(layerCounter[0]), .ZN(n_0_0_76));
   INV_X1 i_0_0_858 (.A(layerCounter[1]), .ZN(n_0_0_85));
   INV_X1 i_0_0_859 (.A(layerCounter[2]), .ZN(n_0_0_86));
   INV_X1 i_0_0_860 (.A(poolingCounter[0]), .ZN(n_0_0_259));
   INV_X1 i_0_0_861 (.A(poolingCounter[1]), .ZN(n_0_0_279));
   INV_X1 i_0_0_862 (.A(poolingWindowX[3]), .ZN(n_0_0_393));
   INV_X1 i_0_0_863 (.A(poolingWindowY[3]), .ZN(n_0_0_395));
   INV_X1 i_0_0_865 (.A(convWindowX[4]), .ZN(n_0_0_396));
   INV_X1 i_0_0_0 (.A(n_0_0_428), .ZN(n_0_0_397));
   INV_X1 i_0_0_1 (.A(n_0_0_278), .ZN(n_0_0_429));
   MUX2_X1 i_0_1_0 (.A(DMA_filter_number[2]), .B(n_0_570), .S(n_0_573), .Z(
      n_0_576));
   MUX2_X1 i_0_1_1 (.A(DMA_filter_number[6]), .B(n_0_571), .S(n_0_573), .Z(
      n_0_575));
   MUX2_X1 i_0_1_2 (.A(DMA_filter_number[10]), .B(n_0_572), .S(n_0_573), 
      .Z(n_0_574));
   MUX2_X1 i_0_2_0 (.A(DMA_read_write_filter_bias[0]), .B(n_0_567), .S(n_0_569), 
      .Z(n_0_578));
   MUX2_X1 i_0_2_1 (.A(DMA_read_write_filter_bias[1]), .B(n_0_568), .S(n_0_569), 
      .Z(n_0_577));
   MUX2_X1 finishCNN_reg_enable_mux_0 (.A(finish), .B(n_0_549), .S(n_0_560), 
      .Z(n_0_579));
   MUX2_X1 DMA_start_reg_enable_mux_0 (.A(DMA_start), .B(n_0_550), .S(n_0_559), 
      .Z(n_0_580));
   MUX2_X1 i_0_3_0 (.A(poolingState[0]), .B(n_0_551), .S(n_0_553), .Z(n_0_633));
   MUX2_X1 i_0_3_1 (.A(poolingState[1]), .B(n_0_552), .S(n_0_553), .Z(n_0_582));
   MUX2_X1 i_0_4_0 (.A(convResetState[0]), .B(n_0_554), .S(n_0_556), .Z(n_0_636));
   MUX2_X1 i_0_4_1 (.A(convResetState[1]), .B(n_0_555), .S(n_0_556), .Z(n_0_634));
   MUX2_X1 convState_reg_enable_mux_0 (.A(convState), .B(n_0_557), .S(n_0_558), 
      .Z(n_0_637));
   MUX2_X1 poolingReset_reg_enable_mux_0 (.A(poolingReset), .B(n_0_563), 
      .S(n_0_564), .Z(n_0_643));
   MUX2_X1 writeReset_reg_enable_mux_0 (.A(writeReset), .B(n_0_565), .S(n_0_566), 
      .Z(n_0_647));
   MUX2_X1 convReset_reg_enable_mux_0 (.A(convReset), .B(n_0_561), .S(n_0_562), 
      .Z(n_0_648));
endmodule

module main(start, reset, finish, clk);
   input start;
   input reset;
   output finish;
   input clk;

   wire [15:0]DMA_filter_number;
   wire [1:0]DMA_read_write_filter_bias;
   wire [15:0]DMA_start_address;
   wire DMA_start;

   RAM RAM1 (.enable(), .clk(clk), .address(), .write(), .\output_data[0][0] (), 
      .\output_data[0][1] (), .\output_data[0][2] (), .\output_data[0][3] (), 
      .\output_data[0][4] (), .\output_data[1][0] (), .\output_data[1][1] (), 
      .\output_data[1][2] (), .\output_data[1][3] (), .\output_data[1][4] (), 
      .\output_data[2][0] (), .\output_data[2][1] (), .\output_data[2][2] (), 
      .\output_data[2][3] (), .\output_data[2][4] (), .\output_data[3][0] (), 
      .\output_data[3][1] (), .\output_data[3][2] (), .\output_data[3][3] (), 
      .\output_data[3][4] (), .\output_data[4][0] (), .\output_data[4][1] (), 
      .\output_data[4][2] (), .\output_data[4][3] (), .\output_data[4][4] (), 
      .offset(), .input_data(), .finish());
   DMA DMA1 (.start(DMA_start), .reset(), .finish_read(), .clk(clk), .address(
      DMA_start_address), .offset(), .read_write_filter_bias(
      DMA_read_write_filter_bias), .filter_number({uc_0, uc_1, uc_2, uc_3, uc_4, 
      DMA_filter_number[10], uc_5, uc_6, uc_7, DMA_filter_number[6], uc_8, uc_9, 
      uc_10, DMA_filter_number[2], uc_11, uc_12}), .\CNN_output_data[0][0] (), 
      .\CNN_output_data[0][1] (), .\CNN_output_data[0][2] (), 
      .\CNN_output_data[0][3] (), .\CNN_output_data[0][4] (), 
      .\CNN_output_data[1][0] (), .\CNN_output_data[1][1] (), 
      .\CNN_output_data[1][2] (), .\CNN_output_data[1][3] (), 
      .\CNN_output_data[1][4] (), .\CNN_output_data[2][0] (), 
      .\CNN_output_data[2][1] (), .\CNN_output_data[2][2] (), 
      .\CNN_output_data[2][3] (), .\CNN_output_data[2][4] (), 
      .\CNN_output_data[3][0] (), .\CNN_output_data[3][1] (), 
      .\CNN_output_data[3][2] (), .\CNN_output_data[3][3] (), 
      .\CNN_output_data[3][4] (), .\CNN_output_data[4][0] (), 
      .\CNN_output_data[4][1] (), .\CNN_output_data[4][2] (), 
      .\CNN_output_data[4][3] (), .\CNN_output_data[4][4] (), .CNN_input_data(), 
      .RAM_address(), .RAM_offset(), .RAM_write(), .RAM_output_data(), 
      .\RAM_input_data[0][0] (), .\RAM_input_data[0][1] (), 
      .\RAM_input_data[0][2] (), .\RAM_input_data[0][3] (), 
      .\RAM_input_data[0][4] (), .\RAM_input_data[1][0] (), 
      .\RAM_input_data[1][1] (), .\RAM_input_data[1][2] (), 
      .\RAM_input_data[1][3] (), .\RAM_input_data[1][4] (), 
      .\RAM_input_data[2][0] (), .\RAM_input_data[2][1] (), 
      .\RAM_input_data[2][2] (), .\RAM_input_data[2][3] (), 
      .\RAM_input_data[2][4] (), .\RAM_input_data[3][0] (), 
      .\RAM_input_data[3][1] (), .\RAM_input_data[3][2] (), 
      .\RAM_input_data[3][3] (), .\RAM_input_data[3][4] (), 
      .\RAM_input_data[4][0] (), .\RAM_input_data[4][1] (), 
      .\RAM_input_data[4][2] (), .\RAM_input_data[4][3] (), 
      .\RAM_input_data[4][4] (), .RAM_finish(), .RAM_enable(), .FB_write(), 
      .\FB_filter[0][0] (), .\FB_filter[0][1] (), .\FB_filter[0][2] (), 
      .\FB_filter[0][3] (), .\FB_filter[0][4] (), .\FB_filter[1][0] (), 
      .\FB_filter[1][1] (), .\FB_filter[1][2] (), .\FB_filter[1][3] (), 
      .\FB_filter[1][4] (), .\FB_filter[2][0] (), .\FB_filter[2][1] (), 
      .\FB_filter[2][2] (), .\FB_filter[2][3] (), .\FB_filter[2][4] (), 
      .\FB_filter[3][0] (), .\FB_filter[3][1] (), .\FB_filter[3][2] (), 
      .\FB_filter[3][3] (), .\FB_filter[3][4] (), .\FB_filter[4][0] (), 
      .\FB_filter[4][1] (), .\FB_filter[4][2] (), .\FB_filter[4][3] (), 
      .\FB_filter[4][4] (), .FB_index_filter(), .\FB_bias[0] (), .\FB_bias[1] (), 
      .\FB_bias[2] (), .\FB_bias[3] (), .\FB_bias[4] (), .\FB_bias[5] (), 
      .\FB_bias[6] (), .\FB_bias[7] (), .\FB_bias[8] (), .\FB_bias[9] (), 
      .\FB_bias[10] (), .\FB_bias[11] (), .\FB_bias[12] (), .\FB_bias[13] (), 
      .\FB_bias[14] (), .\FB_bias[15] (), .\FB_bias[16] (), .\FB_bias[17] (), 
      .\FB_bias[18] (), .\FB_bias[19] (), .\FB_bias[20] (), .\FB_bias[21] (), 
      .\FB_bias[22] (), .\FB_bias[23] (), .\FB_bias[24] (), .\FB_bias[25] (), 
      .\FB_bias[26] (), .\FB_bias[27] (), .\FB_bias[28] (), .\FB_bias[29] (), 
      .\FB_bias[30] (), .\FB_bias[31] (), .\FB_bias[32] (), .\FB_bias[33] (), 
      .\FB_bias[34] (), .\FB_bias[35] (), .\FB_bias[36] (), .\FB_bias[37] (), 
      .\FB_bias[38] (), .\FB_bias[39] (), .\FB_bias[40] (), .\FB_bias[41] (), 
      .\FB_bias[42] (), .\FB_bias[43] (), .\FB_bias[44] (), .\FB_bias[45] (), 
      .\FB_bias[46] (), .\FB_bias[47] (), .\FB_bias[48] (), .\FB_bias[49] (), 
      .\FB_bias[50] (), .\FB_bias[51] (), .\FB_bias[52] (), .\FB_bias[53] (), 
      .\FB_bias[54] (), .\FB_bias[55] (), .\FB_bias[56] (), .\FB_bias[57] (), 
      .\FB_bias[58] (), .\FB_bias[59] (), .\FB_bias[60] (), .\FB_bias[61] (), 
      .\FB_bias[62] (), .\FB_bias[63] (), .\FB_bias[64] (), .\FB_bias[65] (), 
      .\FB_bias[66] (), .\FB_bias[67] (), .\FB_bias[68] (), .\FB_bias[69] (), 
      .\FB_bias[70] (), .\FB_bias[71] (), .\FB_bias[72] (), .\FB_bias[73] (), 
      .\FB_bias[74] (), .\FB_bias[75] (), .\FB_bias[76] (), .\FB_bias[77] (), 
      .\FB_bias[78] (), .\FB_bias[79] (), .\FB_bias[80] (), .\FB_bias[81] (), 
      .\FB_bias[82] (), .\FB_bias[83] (), .\FB_bias[84] (), .\FB_bias[85] (), 
      .\FB_bias[86] (), .\FB_bias[87] (), .\FB_bias[88] (), .\FB_bias[89] (), 
      .\FB_bias[90] (), .\FB_bias[91] (), .\FB_bias[92] (), .\FB_bias[93] (), 
      .\FB_bias[94] (), .\FB_bias[95] (), .\FB_bias[96] (), .\FB_bias[97] (), 
      .\FB_bias[98] (), .\FB_bias[99] (), .\FB_bias[100] (), .\FB_bias[101] (), 
      .\FB_bias[102] (), .\FB_bias[103] (), .\FB_bias[104] (), .\FB_bias[105] (), 
      .\FB_bias[106] (), .\FB_bias[107] (), .\FB_bias[108] (), .\FB_bias[109] (), 
      .\FB_bias[110] (), .\FB_bias[111] (), .\FB_bias[112] (), .\FB_bias[113] (), 
      .\FB_bias[114] (), .\FB_bias[115] (), .\FB_bias[116] (), .\FB_bias[117] (), 
      .\FB_bias[118] (), .\FB_bias[119] (), .FB_bias_or_filter(), .FB_finish());
   CNN CNN1 (.start(start), .reset(reset), .finish(finish), .clk(clk), 
      .\filter[0][0] (), .\filter[0][1] (), .\filter[0][2] (), .\filter[0][3] (), 
      .\filter[0][4] (), .\filter[1][0] (), .\filter[1][1] (), .\filter[1][2] (), 
      .\filter[1][3] (), .\filter[1][4] (), .\filter[2][0] (), .\filter[2][1] (), 
      .\filter[2][2] (), .\filter[2][3] (), .\filter[2][4] (), .\filter[3][0] (), 
      .\filter[3][1] (), .\filter[3][2] (), .\filter[3][3] (), .\filter[3][4] (), 
      .\filter[4][0] (), .\filter[4][1] (), .\filter[4][2] (), .\filter[4][3] (), 
      .\filter[4][4] (), .FB_index_bias(), .FB_output_bias(), .index_filter(), 
      .DMA_start(DMA_start), .DMA_finish(), .DMA_start_address(DMA_start_address), 
      .DMA_offset(), .DMA_read_write_filter_bias(DMA_read_write_filter_bias), 
      .DMA_filter_number({uc_13, uc_14, uc_15, uc_16, uc_17, 
      DMA_filter_number[10], uc_18, uc_19, uc_20, DMA_filter_number[6], uc_21, 
      uc_22, uc_23, DMA_filter_number[2], uc_24, uc_25}), 
      .\DMA_CNN_output_data[0][0] (), .\DMA_CNN_output_data[0][1] (), 
      .\DMA_CNN_output_data[0][2] (), .\DMA_CNN_output_data[0][3] (), 
      .\DMA_CNN_output_data[0][4] (), .\DMA_CNN_output_data[1][0] (), 
      .\DMA_CNN_output_data[1][1] (), .\DMA_CNN_output_data[1][2] (), 
      .\DMA_CNN_output_data[1][3] (), .\DMA_CNN_output_data[1][4] (), 
      .\DMA_CNN_output_data[2][0] (), .\DMA_CNN_output_data[2][1] (), 
      .\DMA_CNN_output_data[2][2] (), .\DMA_CNN_output_data[2][3] (), 
      .\DMA_CNN_output_data[2][4] (), .\DMA_CNN_output_data[3][0] (), 
      .\DMA_CNN_output_data[3][1] (), .\DMA_CNN_output_data[3][2] (), 
      .\DMA_CNN_output_data[3][3] (), .\DMA_CNN_output_data[3][4] (), 
      .\DMA_CNN_output_data[4][0] (), .\DMA_CNN_output_data[4][1] (), 
      .\DMA_CNN_output_data[4][2] (), .\DMA_CNN_output_data[4][3] (), 
      .\DMA_CNN_output_data[4][4] (), .DMA_CNN_input_data());
endmodule
